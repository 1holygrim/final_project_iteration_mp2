XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��46�̟�k+Z��9�����\؈���ܦjkN�,D>���z���*˲,��䗿A̒:a'��4��z�լ䈽��_Ὁ�ՏP%�E�@dQ��M>�@�n��3��<i��[�P�xj���(��L��{͞Ce���� ��m�y�ӷ�T�����o�沔U��;���b�EJ)�7&�-ًz��eF�q8H�4�@DЈ����Jw�Q��H*����[�,g
��͡�
�b����.j\��>\���aF\�Z�h͐��_�IZB[1�Q�a���)0���W�Ȭ|��F�p�&��ik����1�ЧQMiKyf�I۹�cf�NHP��rJF���>�]���:ٔ5��0~s������ed�
]|�r�kX
��t���������Y'�(�/LqՐ�%q�X%K�yQ~ $
��ӑ��\_^x�V>d88K��`�s$�XB����?�PD}�x���//�7 p�/�g�����-Nu��A\@-��e5���-�B�W�y��ы�6p���7>�����~p���.�)71]���&n�P�;7�R�C��I^�B�ȖF��6v�Ț�����@(��3��H"5.ImzF� jQ7t�j��1��P�V��zS̖���2��O���z}�g�+3w�<�' HH�!�}J����H5���jV��ঌ@���>5�t���/�H#�5حPv���2�5�����{�+�śId<���]��Z��-����`+��9N�jXlxVHYEB    b229    2170�d��pA��̷um.��埻�װM��%Q�}�0��a�UP�<� 6|(E3��K`�V�}�� �GR��=�:��vΎ�i/����l��}�k���5c�+w�^��u_�f�D!����S�>��#�����iI�S��S�W�9&[�f�Y��z�6���d/M��b訠�4��S�'���m�a��6yO
�%����=�gn��hO\�9��_5�R�#��!a�M���"'�p�����y\�T����j�gڙ��=[i���k�Jl�g3���@�e�K5����{ �8�d:�[֩�{o!���a��b?՛�J]���/9/��/������Q�i�5��LZu�]��4ѷ�'�Y�N���/:�l�Wl�-G0Q��́�HP�l�گ�w� R�J�\�nz�޽M��")���2Enssa9t����$A�9@��)L">�F�k"��6f�L#���\���9�"��LIP;ޜ�%|�=�A{7�p�&���*/�(�c�v�5��}�2b�I@ߚ;�vSTh��$�1�����G�!hIJ��6�r�N���&^�**W���X�1Z���)ޥ��#��B��dӗ%ӧS�Dޯa�1�i�����w��Y����. �(��6���G�����O���;N�����G��'�!�t*�6ɑ���W»[�$���������\�7d��,�'E<)�QgXߞ=��gHcӎ�za��ӼZ(-�,��#��7O���:|�ګr0X����Â!��������A%z�o_��oR2�W����K�ҩ��P�b��(�4����r�߭��4�̳VN���hy���v�y�p��_9(>+�O �E��I����\3"lf����GR�;��%9�fԑ~N�"�bE���TL��4ԒW�0��!�E���^M��D#pj�HR����,����gR;�Ad��h1I�����>{mb�Ơ������s'���� L��o��9����N��_��g�Kڕ[`��TK��b��<�1��l��<���BH����2g<hKR��lV�/pQ��$uutb;R' }8�u��޺*� \���x^hd����11`)�uB�n�[�4.�i5
���
�Y Fǟ�_ry���8�[z ����DdMb86�>;D��u�m����IS�e���Ɩ��*���Xq�v�~G�̊
h
���PԵc��ɮ��r�a �5��F�H�S'�0�X�rV2#x�5Q��d3,6�_��()�h�-��4Ż�J���F�-�p���2j����)��E���#Z���G�ɤ�w�YY?����:��W��Tw�t|��}�n���@�?�0��t�Tj#���4������w�W`�e��q��Ǉ����uGi�w悯����	�{pZ���k�&:�V�A�T{���ۦ������yn���.��6���l��|+���Tgn�jz��hn^��(kv�j\A����p�+M��jMĮ:��s�����
�|ӣ%��ɝ�0:A��6p'?x�(nW�W)U���C���/�޹���jr
���X4��qk��p��N���r7�D�RU7Ip\,B}g(�\��Mt�]V|:�XsA�9F��֤��~� ��yc��,�͕5�QW �ӏ��_�v1��EGO�du2˄=����8�#<�e�� ����\�0�NVC���m���?��ԑ�r!��>�9�p����@<�1��.�5��hq������`L�w�X�6"�Hu�-�u�lq�M�'6�T�$%�:����]�12����de�pt^���*���|�OܾV�ʙ��Yj�υlQ��+�# �Yp$h,8��%U�;6��/=@$�$8ӹ�)(ۭ��ܫ\�t�VԠcWZCz�L�?GK�3�e�T�Y��?�� �G��W��G�[0�1�����/܂�@{~�b�E��-<�J�h�45%���1}~҄�+߯�x���͔u�Z"�3��%�������b�t�z11?(��0�=�En�S�ר\p�INc�	y�Fg�r�^m�R���.'p�v&�[�Jͻ�āS\�{Gӏ�{JɩY�����k��(�P�@�N��}�i�����{م��Ў�;��O���Ƣ���L\̘X��էl� ������fJ������x�s�����.<���!A!�ul����`�*ִ��7��/�/��bʳ�nN�[V��/�Dfn�!�}Wsh������	p�Y��CS�^k�<�zp��4-��w#�Բ��u]��J�������-��Ǖr�2��X�C����NhK���&\��$�4��ɾ�q_/�o�=qgا���O$(���2)��I�e #���mzk��$צ�v�n�BZ����P-��@�Y%P�-����4R1�
�kV@<���6�rڙ�gó##�#ݧ����Y�vb��+�����折��;����0�u�����e���a�,S{r�2��PΛ�p��<C����%��Į�zE�)
*t��:bH��j���D=��֜���V�u�8�_���%���J�]�K�81�4Hꭲt/�p��G�X):|�(�dlܙ3Jʒ�s50�8^l��kaP+��5��YW�RI4z��>�Ivh��B�V"B��[	�f8�� _�8I&�U��g����ev�gA���3����b6b�SQF��y�ͱ������Ů���~#Kg�}�÷X},�k�ć�|�*����&��}M���W��(�f�`B��hX==dp���_�{i�A�/Jw�����������ұ��~�b�c�M����y>��������g� �d��R�F�M!�a_��gJ�:=ו��Dp8���R�6}��"�4���7�?����U����z#?�ц��t�W�um�h��I1�jBC����2-�*��@[��~�׀�����$����Ϥ������l���6ttA��@�B��Pk!��\w�Q���5`���r������\0'uv�qVB\��+��)�=�[2��9@����U�%�d�j֍����)�j�y}���\�1�/���r��{}�Yۏ�'���szZe)�6C⥣��na���.L|�ڂV y"�0��Nn�`�ܘ���p��/��S�*�z²�)IX���1(�P�$*;����M�򪤯��U�o����8��dVD@d��a�)&C�QR�!���m^��� ���`+��S�:���%#g/r+,(.���`��e7�!�Yr��a�=�1s�}�{H"Z�N�VB�+�Y�:�Sf��2���ԑ��)e>.v}�ϱ�҂�ţ��$��h��ۧq�����z������l@�+����P 떸?�_T3�y.��R;�z���#^�*!�*��zg��P��s�c�P8�JG��{X�m!���g�:�%1�F���!եV4����IeT����4��N_�@��V���OU]����B�X����꾟���[��P�H��\����#ov��й1WZ�b�� ��Xh���#G�ށ�5۬?�Ug6*`��l���A���$����$5�������qU!��.A`�5���*�mA���� �R�7��f��
�5��j��(3��K���p9e�ݼLI\��z�{WIwy��y���pL�&UJG������@��r�m��EF+5���S��3�Cw��1j®ZX5�.o��1e���za,rJB&꟎��>�/�\�����1h��Iݯ^�mͅ7Vʁ�[0��s@�U�����S��t��BA	�D?��]� ���#vFF0ջ�w�����
��}
0�݈\)hcߚU��� ̡�ZW�����%��o���?�j0Ea�%��R�z8�����ة��\`t��gվ�:��#��i.���i\�p�?�t���Z���O|(Ƶ� ����3;�ۆ#�{z��	��{r�?l�h��kN_68�e��a��fǑ`s#\1;@�*Ll��/�!* 5��Wi���̅�F�[�w������J;�Q[�>ci�F��/�E'r�9\%��!~���@k}<���D ��X�� )S�)h�h��V��%!K��&�a��3���X��W��$:l�|H�
�茅2h	_Q ���/�0��?�*F���6ί-�drn|~�6��\�IP04k�gd�f��E���U?���G��Y�ݱ"��1pw�I����A �8�k�g��W� ��3�3v9�U1|-i=�ws�E{���s�O�U����D�4�hڑyw�V�~	�oun�?bW°m�Iw�$���2����H獠G��c�*N�!T��b*��PR���?}!-�������a9C�R�3�6	��f��o�6������s�س�����/�?:M�S�עL���3���}IN[X�
/M�Q~�6iTq������� �ՎS������!���'"��%u���F~���%P��DQ�y b �^�y�<P���&�q�^�J��8�=0�չ��M���Dr���:BQ�}�O�����e���`���LO��!�C�\�Ȉc�]�.�!�4/��+q'�M�1��җ���[�k�`�����[�Ƕ� ���P�����Dn��t��H�XV���c�,mن�Py2�&�_p���_z,��kK�f�ֵ2�J�Y��U��HK��֐�SH<��gm�j>"���ʘ�'�).��T��D��c J8�3<^s��8v2ů�ٙ��F��U"��=�fD,:�l�q��H�l�������$_)�ģ��~�����A�[�4z�2�g��aR%��r$8�:kHujK�?u#�*Ӯ7e��G��,֭&|:�V=9��1��q��?
hrlj����\i�1���Rgۈz�\��רd"R��EW<��Eq��zܼG{�m��,���4�m�t�p��\�������]r:��׍���%6Rs>:�.^H_%��U^��d�4YY�X�D?=V���q1���<Tq���{�7YQ?1oJW��Y0B����o�7ᬮ��j�����q3"�h�k~����[�L$5��J����l�~�l�[�%��?���)�֤�ĸ����Đփs�a4����b�{\����`�wUPf��o-���A����-�j��+ ~�a0m9w�hO�����N�ہ:ӄWkO���4*�j�p��!�գn���q.�`�;�%d?dAK4�~6S���AA����"[Z�����íH�~i�]�؊��lQ��%˻3Y�b���X=ѕ�[�V��`�W՜��� ݶ f�v�F,�+U��v��fU��&k�:��fq�Y5�x���n��k^հ�B�L�����ꮷ�࿵dgI��7�|���*ܿ�%��9"�$Rc?�T!̟7N��:�;Q�w1�G/�Y/�@�"e�ڸ!�42,��2�p;�f�����'l�+�ܩ�$��qNq�!�AW=f��ϖ{\Sjw5-���	��n�{�)�^�#pԵ$�
n�Ϳ�R���9i[l�&.Vb*"��D�q�H��NDi��`�=\֘!I�!������TO?��=a�n��C���9T�����\_���tО��}������q�S��8�8��sq;�.w�\�$خ�tX���+ ��z��!��Q�W��q�lH)q� ����?@�B4[�z�#���D�|�UE"�(BW��Ws�I�Yn�4�ŉ�v򞪤���j��Q�\�Iſ�����jz3� ���ڄ��� ��Mɨ������n4�~PC��	ڥ���0�rΒ�����wJ�!{¨u�L�"]��v~���w��1�~;I-؎��Qp�e�4����κ���V?�~vc�K��Fyee�<�N&�(pꭢd���p�;~P@��ɔ��z�X��p4��YSQ��15��3�-����S�����o�7��xG������jxl�:�(D���L�=; d���_����A�=�n9�$9g����N�v5��
���|DUW�?�"��b#�K��k��Ĵ�BS�徙��-��хc )&y]�bJM�ռ��w[�Z�j�Ia���ѾҎ�Q}�wǷF�nR8���V�@�A�gi.�j��i��y��ɑ})�=J����+��c'�ns���E� �W{|�o�!_��G��q�j���ڽ�!8d|w�.B{~l\����wb�8��Y���jJ�K����ur9nO�-ncs[׸�8c�	�^���7�(��I�
�'��*��U�ǌ��]X�7O1x-"cǆ�:u��c4��6����M����lA�� >�B*l�*���з_X���do-E$�8M+�/�`����ڏK��4��W�_LO,E8�#����1I-���Ֆ�O@�
�}�,4]���e��JzOb�%F�A�hN>}D;W����a��?٥���L�|������?�7�PL�� Ηd���~Sw��Z-����W�(��^��d�_��uN����!�����w�m�/�,���l�!�pӫ�{{� e�]>|����,mٖ������˃Ck�:�dƄEG<�E�YS�EI�蓓잩���� p�7$$�p��}g}�@��r�h�
7����&�2
+ɬ*�A�J��~z����E�H�\�M�x��K��3����	����	�������S�ʧYHu13��xQ���-�E���MƏ2�^�R����(�{}�p/��o�I� �(&2��.N�ո�i��_���S�ϴ�azqNZ���f;���[8��GqP�X�\�Vgne�dV�{Y���ۖ� �� �Å%�����s�a��4���5يx�)@<9�~U�[��3�"��W:(�z"@��ng���n�%�ȱL.|���C$�sէ��YUL�0s~��@>w�
j�v8pR,8�1ޭ��c~�V�xjCX���6��lP��,E#ȃ���-���O2�*L�o�l������)� �R�� Z�}��E�9XD�"�[���A;CRx�f�(_�1VRg�-F��Kq�I8Ae({�м����"�
������j���DW)���G`�% N-����L���c��&�#������B��v����.��k�p�-��6�@�K�e��Ā8X���X�y������i~j]<���Y��j�+}tI=p��t�SK`�)q���ʾCV,�ZUFm�š�ƨçP��O^=�j��~�7���I�|�j.�I.d���g�ۨ�vG�7W��v���F	�nb����좱�<�3���DH_4����YP����)쬽�p��ͺ�lֻ�T�AT�~u�OO\�z�h|=sV!�>���<OK�v�)�bȧ��߼�5ޗ4��?3��� W 0c��0&q��z/م�VU�B"�rb{�@�Z������Op	o�Eܑ
�0�V_\f@(}����w
�Yr��+/�|oL�\��F�U:���I���C�������v���s��Zv �U���ܰ2&<��Ӓ�5����W��-�y[=@u#<x���#��me< ~#."�VPr�D-���8��^'��m�j}{�&���,�:C�b�G��5A`�H�|��ֳ���-�xK�B��޿��I�d��"@���Èa�z����v=�5O�(�qW{N����8� �X���4��[����z���g��$z�	�)���c�d���Ҫ^�x%���0?�6W�bDr���!��_�����.&(��x�}�O���Pww�+y&)��Y���x<���!h�_�j��(r��iXY�J�H��Ko���p��O_�q��ŏ��5��� �5�r���9���ygwc�	�\-� �S5	l۠1!�vy�R_��#A��R������9+I�k�E�����=���~�� �c���������*��;m�tX�O���_����?lQ�j�`,��n��3��[@'Y�WQ\�BS,mFmc��J�V�%/*�����ױ���0�/L�8��g�K�+c���Y|5�&��B�Fh3|	��iU������"c�Y�����M��	��C�{A����`����^�"V&zC9#�жD����߮�	��Q%VkStZ�qƦt��\��vW�
�w[µ���M/������<��֕đ�v�;o��=����CGڌ�>R�q	Ѫ������E���\�/�E�J�Ω�8�P!���0��/���*&� K̋ .ӭż�s��vFϜu��9O�7�C�{qZⵅ��Q�]�_{f�&����g���v&�/<�RݮBNN�d�����80�.��D��K�ˤ��t���x�47���k�=���65���7�i��%�n ����R��G�M�j.�I����_3��4�����o�@)3\݋�i|G۽��1��DYM[Xm��^NP!����