XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���g�s2������5�H��Yi��\X-xi�!/y-�WD��l����d��
�����#��8-������t��tA�LA���Ɠ����>�y(�dr���Ȥ4["��B����֚�o�M�6�n��ݣ�;���Y�~psv��Q��q�̃��.�h�ub�8og�%Z6�ܬy�xmX#"��OGS��T�R�}��k$Bh0؄��ΟA-����t����(���Ϝ&NgH��ӹ��UI��X��/��L�)`)����0�^�1XCMʧ�aUUI�aYzc~�?�$L�Њ#���#��y�H�E�5�~�_"{�R+[%*uY�=��ɩF��Ш.Gi�c�<��#sA"e顱�F�A��I��9!��h� ����U�1�߶��J^�0��i��tS�+�5�v�ld�D�%�����.�^a0 &�����Q ���mm��_r/4�M�'�������d ������{�QwTuDP��i�{�BO��b�#�7>MB���=W���Ȟh+/}ض��7
u��c;���Oj倌���7qO��n;��a3�yp�ļv���T9���ʨ#T)D����<wԥ���P��[t�%��Pf:���h�.%��#8b���Q\9H��A���b�`��uƏO�]	�{
A��Ⱊ�sQ�.��)��:��-�i��3Pye�;�[,o��$?5�m0�;S1:�Uq�mߐ�Msĭ�ٙF��t^��ٟ}����,��8�.�iML��)XlxVHYEB    95d3    18d0�����(����k0^AI��DQ�F�	�8@?	[�.S�~ݻ!ڻ����eDց��D��5�^i��o�=ر�k�`��=0e����4�m�H>	�yD_�)�k�o����~
�z��FE�:�H|�z�(�&�ƺ`�n��(�b��_�[��b��y�Vg���g[�J��_�h2Z����o]i�斿�z7�ͩ���ZF���Y�s��j����7^kmDg�v���/� �x�.��s�p�mdpD)?]]�g�Dj��	0�����S
v�;E;�>�rڶ�T�sCN0�N�a��b������'�A�.�n� �Y�@�X��w����q��yN��Q�Y$ �w�)bh�;���k'�L�����)�˿>"�&��7�T��<�BT�{`�3!����!��|��Aڍ�[;r,��Q�ܔ�M��_]�NL�7)�,`3j�B'#�qwf5�����.ʍPp��*5�RvW�������v&<1���
7ߦG�7�v��%h�Cl}�i5�u
cA�f)O͕��qIS
��$u�iR&|���Xx��d�vU٭�^�a�V�2ه9����]z�SM�~�� �,Q�hȄ������v�l��Mf ���.xA�rpRC���Vʻ
HA���s%|�x���0$kMH۔�ow���*��IT��V��߃kc#�w_�
9p�<�E܌����2|����؀�P���4�H~�ǉE��6
e0/��6�}2?�G5焷���̦ꝩ�������U��mb��-6
/��1߆3��(�zC
�K���~g$�d��A�'P����Z!��4�H��S�s������<�w���$Ao,-�N_$�D^�������f�Fy�a�sf�e]�]�8fM�RE�OY��c�xW
d�K��:������AH�HSt��A.����öp��DƬ�׊�7���K�cq�+��e�z� Xm�l�C��dz[d��:a�U��#R�e��Q��E.U�I��G���r��" t�E��~�8�"�n�c�.��KQ���?��C��ff��(�'v�D�kDJ�f�W�b��gh���*{*Ѹh&�����_?ƾ4����@��.�P��9�eȿ�53l���m ��>�5��E��	ْO���R���:��g�����lb���Y���&C��+�P���Ħ���9w�˓��C���2��S.�	Y�V��1��P�r4�t����h9}�V� �7��
�2]��9�-39�ŷ��I�4p
�͜X�&��j���䖁�H��H�vԈS��A~�h�>'T��[��`���Й��.���͂�.�������J%p!�w���J`U?�ɴ*�C�|Nc��qLQ0Tәd��<������_��+�rkg9��|��(��$ =�|�{ �@ n��I��:��;?z?]�ո*H��p�uN�y��t�p�0eՍ4�1d�WP�6â��xm&/������v%��",�q+^�2�;b�M�݄�%�HbD�n�����9N���s��2�.-i=��v�
}�+�#
7�{��ix��Sd��']�ޢ���@�� s�D���7U]�iE ��S���+M-k��B)��:�u	� ٤�E��|�ޫN�ha�h��.} ڜ'�� ���yHxI�fD�p������Of�smt��f��<[�ߛt�ӕQʩ:!n5*2���y��_!)��^V�r�	�KjgqT�����w	�`���w�%AĲR��L�F 8�R�Ѯ���tM2�99.6�i���&�����)�kQ�$���� �bl�Ï���.\�w�F)�u��fw4{G��D5[#��Y�W�@1���j��(}�� <=�~ݻ��aL�J#�Ю����xM���Oʔ#�ꭅ���(��L��/!ZT\1�QT���� E��;�8�?��C��ۻ³��b����d���!�o���{�L��r���XR�h��O���X+�L6 v�F�Y��jsYY��F��w��63��S�nfT�� ��Z
,1�=��흉��#�F#��[�A�O�^���TY܏���l��"�c��{��ݙ����2�N˽N�|l�O^��a� |<�A=�}V�4�������Ƙ��&�4\W�����mm���ΑJy�+"��v$^	�+׿���{�g���z���po��B�\���+�V8
��c���5�����Ef���
�$� ,���;�9VP��[�}�SQ\\�3��H� �r���>Gl���^�S�f��D喆�Θ=z���j���N'(p���K���n�q	��V�K�J�T1�3��#)��ΐq�7ܨ�Lґ�E�_�1��S�b��U�<���/��Ygӣ�V�������j H���]{
��;.�A���uЧS�O�o���	�ͱ���q�|3��O��!�68�̚A<!��{��l�e;�48�(pŜ�����c𗁘�=�`�|��mD�!s��5����(?�v��:�vʄ��(��s�H (��po�=f:�t�b�w�"4\�֎r����_V�����ߢD��nQcg�v)�]��k��-�77>CA�����S���cA�\_�<jQ2"���䓩Z����uZ�0��&�$�~�w^֚�)����N~���)*Y&~�J��n�ŵ'�D`Eaү�4�������r�f��]n�F���/W��kuф�.q]i�f�di� ��)(�~�ŕ��TlSZ�q �d����_퉈K�2MHFD�A)�̰7;{K�����Y^��p��Q˦���U\�BQ�t�f�Jmv>ߑ��4A������wp��U4.]D�-�(x��$SK���Vz�>Xh�ܮ��.��͘���W�����*��=��5��or @��3O����Xk"{o���7�0�y�f�q�.͘&�/@㋎�v:�2�m�/3�`���E���5�Β�W>�� (�1����o���>����/��xu��?��Q)�c-�h��w�pl{�q7p0�u�$lo_�ү��!�LΉ�5IB���}4��?��`�\�9��Jۤ�����Y*��a�h�=؃n5�|�ƶܸ�����R�.+��+����x;�S?��=��|$�m�#������ê���7���}� ���L!������9�z߳���i'�ų{i���՞\��/�F�o(&�RУ^�!�M��ӏf�̚��G}|�&c'G�;�_�g�%���k��E��qU���2����I ��0��+�h�W͠�G>�N�u�7�6sF	�پ�Ņ_���]��&���r�x�=[�٧(3(x&�Y<��a����	R@�f>L����3�qw�;��
Q��=o��v�G��A�L���R3��4e������4��m2v�E�V�2���`ٻ��4�%b�C)��G���Wy�uޚ�U��Y4
sh`VD��E�MN堃�Q������ʑ�}Z	�	]��BdcZ�`~Jgp��/���c�{FfAQ&�'=�� �_��}�?��z䗼�%#�R���땃�r��[�Fi�A��ϒ|��Œ����E�(T�=�~�.�3�n��[]��&�d�/�wD_|Ǭ��bh�:rbz6i��nj�줿����u�;-?s���C`C��I�-�����*��.)o [j��5��[���l΋�d��G�j�Ga�%jl������	�rOnX0>'/i#h5��q>�[]���(o�f�1�[�u���\�k�P��˦�����=�B�WĢ�ijW,�S�����`�v$y>�$���T8�����\�m�s3H��bOJ�2Μ�$G�ܺ��^m
l!\1�I{ү辱<M��G[TXʎ<������Er�����V���鑹�	�:0u�e"r	fj^;�%3�gءd�(��S!�`�b�#�,�E}O0�,�=�g�~"$����J�$����~�9x0�a���Hw�՜�#2t�o X���'v�vh�1j ��M�@*���a��� ���������>X鿔��t�H �j��bB���� 
�����˅wƨ0+���c����k��s����%gYٺ"ы��4� JMP�J��n��g�K�ה
�ce���(-��������ܖ2�Q��]_K"�@�=��GM�ÿB��D��V!%1k��g���ǰ9���i��ux�QAEu��l!���	��5�99�i}����W�t�^MSoq�`����i"��@7�����T�KXy�s�L�+_�y�
������1=�g!��S5�C�e���������zop�l�TS>�(���͆��*f�pu���󧹩�0F$�&~P��6�N]����Ӑ89����]�>��Ob�l?!���bMsm�(������~賧JN>y	c[&���R���c��2�.b�x���g��}�6�p�MK3&�� PCd�6�1۵��r��v<���X�T������s�Z����e  ��m��j���� �q���8��n�G�](�ai��߶�t��hIZ�?񖕅%�X�5D,p(Y�Q��<*(4���&a�'�W����In���W��9t7E#]l֟vw0 �r��?�	<� #1kSl_��cs��B��B��o�?	ک�h���PL�ۄ#zz�ՒL�r�3&��ɬ���e~�}(n-���sq�QL��i��5���$w�B�m��r�3���Q����{�x�Lx=����R'$u+��L4�$��a�Jp�%��il�c�����f���CQ[p�x�󛺆/s���dc�<����ì�|w�kU�_�ꄍt�Ce�G��5:V R��זV[]
?�0nI�"�����&a��9LTm���f�)��!wb�&�$<�^�a�'!17U'���m0Q�_�\��i Cwf�10;��11r,I�k�B��9�:�m/����ߌ򳇜#S��{�V"�xn���"��po�#�%�d�0<ư�ЎG�Rs�DoIѰ^*v��ۣJ�ѓ��pթ�?<tw$e��5�,G��B�k��p��ǝ25���,�D�Ezx�I��\�zĸ�?�v�[�䍌*��v�S�Xo��;,*n0�<�7���@VX�e<�K=6[�Ctvc^����"*7�F�Tj^|���E�W�X"	]��z!���;�����M"a�����:�:�Q%�� ��ah㼗�[W���(�]L��c3�=H� �� z��-au��1~�b1���[�KŞ7�/��:�I1�hx�4Ѿ2�~�;�8Q-��&�<R]-�]����#B��8H��h횸ے���5
Wz�s�P�8G$ϐ8�)�j��ڨ���%�J{�T7�dHJI��E�L~��ַ�x6"�$��e���t�m?��q[�b���U���7�v��S�r+�8�~Tz��~�b_�|��y|NI٣�Pj��˙�2��`Z�q~1�CSd�T=�q	�+��#��H��Q��'�2VU,�Z6��;w����2|��D�#��!���"n�]_Uq�Ѩ.{h�O32{,R[�
�/L�;����
�#�x��@6���i����2��\��u����s��o ̇�O$���\V�V�
LT*<�@<���1%��V�p��:��p.�Đr���$�G0�n��$�Y7/Q�jK����j
L�l-z,�����-*4�������0�P�;HQ
y__�K��a���9��r������_k�=����c�<���iL�&�`�jf$�3��Yi��q��mP�.r>�q<u��ˁbv��l��b����ŕz-0�`n�`l���h��xBjIT�
����A�}\���3���$�8�Ԁ�s��d�	����;��4�t񨚄C�Y����W1ԉ�)�<ԭY'�)�V��7�'�W����@��E�K�oc�Yv���=1��h$'�'�0z�v~��~�2w\�h���ӲB���V��&$�EX�"sH�7�{�*�&d�s0�]��B�����.���S�?�7������Z��+��ϻ�`�{���qu֔GI��Ӳ/�������J 10��_�t䤁S���>�W�(�'��+���B�Q;?��Xq�?��ݴ��.�:g��ABuA�I�r�ƍ$ܽ�;4��W=ے���M t���G�[���T����>�I:���9�b�6�Mվ����Vޢ��xK?'��G���ti�q;���2*��;B��E�{��,����ӮD�)�%ٛ�O9�N�Ꮵ���N�����ٯ��Q�