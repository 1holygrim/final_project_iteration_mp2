XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���-F�X�2����Ӄ!`7��sN�L��sZ��pG�w�^���D��7��`ɳE>d����_+����ä=i�;�&=�s<`8O:�c7����We>��p+W8�v�]lٲ^*�[�'|0Zl�3�?�||��	D'���<�����X�`7�,C�h��,n��������6z�<"�*y"��,wگoocF�FS� )hj��[���
S�W�L��d��z����b�f"4Z^6UU	�Iv� ���vn��
�pa�Wd��~Dg]�A��@K�S��!oJ�>:7�+K�' ��u9IZ�����U�hU5Nl��#��T��H��A�}�|G��w�p�
:W2-3���1F�}\������2�
؍<�����ި���"��M�w��a+j�P�ťe�W4�"M�8�S*��c���M�y;8��"S&�찏m�K��v�c81vu*T�=B~�kV� ?bU���\EW�(�@� �k!��\;"�$>C�Ra�t���������6�/��銖O��93�2�XB,)u���S�t[����r���<�q�~Ī�m E!�j��$-"����� ����'T��h�qQR;���$K���������Q��ȫs��Hy�����1��D/wǁ|�}+�����f�eM�u�A��Q��+ k�{����7��͘��u:���G ��[U��i�~�,��J0{�����];�^DR���x=���1pd��J����j�z��G���'��؆j��cLXlxVHYEB    fa00    23d0Nb���P��)�K}�]�����</:&S�����c�O��{�_������OF`�Yo��Z"H{\��������d��fcV��M�9t�K�)�HФ?G�O��� Y�+�5�i	��G]!�g�/q��5�z`�Y'�5�sq�H'Y.UU�t�FDT�2و3�/f�N:�Ї�_n�uM�9�+x�8�2I�qƒ!gjʉ��'e����|`�x�-��9�ܬ�@"�z�'G����5h�w&�"�����V
�GE�ߪ��Km"A4��J�Kg�CC7�vر\)RG��z�e�|��ͨ��A���b�x'������� g��),�8�8T
o���"��+*c)���kx���T��X��9���ܚ�{�>O|)��e��wr��f.��Dd�,̧��Y>Z�����#���ŎN�.x0c��Ȫ�R ��Xq�J�!��XȊ��j#&�P������]�_�mLm��/�)*=�w+D���vf?,h�8
9$i6ŉ���֔�.�%����i��E$;�*D�qP��Ll#�\�0�M��Jw@��X|sP���Nwn�����=��B�}�}��mF�Q��3Yq#̓v�Q��҂p���=k6�_�ז�Bz���'i�D��\-�:�����)�X��}�r{�UH,���Гx!M������t>�go`P�z�NS��ӷq���."w��wx9��,F��p��i��_��%�EE4w�
�,f�N�2̲��ȇ��(a�������fy�H������ ���dգ���yiMEPwl-�Oʌ>�ˊ��W��̘S�C8�_$���rtr���LG@i��~�ހfvݷ���h��0�ՂIye�I��C�C�a<�	0NR�pC�?p�\Z���{����@v��^5��;+�"� �l���s�{�?��"9��㍱m�x��eN�v�*��&�M���b�U��1�n��(|����zϧ��uj�a
�{�[cE���F%z���y1/D[$ԾǛ'����u���4!�As~�-wQ2�'�^O���R�����0I5S}����+����.T�I��(�%�ڌ,��5N�F@�[����Ukt��Ki�j�F#ս5�!��{Ԧ�q$w�U�F�����p��N��Ӱױ<v�[��{��G� �d/����GΦN�N�;�##��l��ݹG	A,ɐ�,�{J�^���S��#�0�KE�go�h᪅��
߼X&?^P�}���*��I�{Jw�M��/B��9�`��{�R�+������f+|�5����>?@w�\"|��� ���X5*��
I��$ �'�[)i^���b���1&K��� =p�~4C�o>&���_�?f�������i���oס��
P�����o�a��0���Tf��7��m��S�R�d.��V�ms�����J���"8d�;�R����ho��'楑�N�6����9b�^T�s)�Җ��N㞯�"%��ݥJ@g�z��b!��j������ȃ'�;4h���:��)z�7v�S/��%g
���`>:���{؍XNN\⾊r�fdxb̊
�=¹�l`Z�[��P?)fbi'@m� �_���e��x�_B���X9"�~��:��WS��E �'	j��r7���!FQR.;6pKuk��d��H��s��4O%$�(\N~L�|}V���.�됅4�x� �}Ap"VE�g�̱�s��v�d���k|���*�B5�8�∇��)<�*��̗�_�>n;�i8�i��Y�w��m��¹?��2�Qf��.��.�Ͻ�TKv�f�O�*���Ӟ)����Ϳ�3�v8��B�e�ţ�w^t'-�k����|s�BF�����9����Я��
݁�����=�W��<2�h�G��UɵB4�pOzI��K6�M����SXK��v�ֶ�դ C��Lax�Ԣ2�(!ϟH�U�e�Я���4 h--��S��\��a�dƠ�W�!�C������"�e����U���u���nx:8��2A8�2�*?�Uzw{6��[��8��_<l����&O���U������,�l�i�er�B��ڃ(�7�{+`����3iL9��~�v�S_�U�J�-X�5ʮ��w]A� -Y t�����������P5�O� ��O%���a�2E%1�T�&ൕ���M��p:2�6��C��u���^�٦�]qZJ�*�0[R�p��[�ҼD�`���0 NJc� ��OB&��.i�Xe�3����`��n�����Z#J`�����mH�EO�U:R�����XZl��*��<R�g]��Srȃ�$�Q��Q�%o��%�E<�2����9h��6% 
S�c��ܗ�/�%��%�����$���"q��p��QH��jvn�Zd�1|}��Ӏ)�����g�����ŴN�O���f�sO_�*}1ƅ����7��9�m���@�<�ο�;x���E�x@�u���XF��b��i�mI�x�ĶwL;���n~�����M����dy`���<�����'�kb����4`�.��2����o�����P"�e�N��r	}�B^N@,�`.<o"χ'�e���6؍�5h��4��z��L������UX��6G�D}��=*�h<�'��Q ���0����6��&Hm�MxɄ羹墨��>P��$���f ��&�q����R�c��<y	����S'z��#��'�+�9��3��;Y/��e�V�gIV���e�~2�G$����(c�/�������r$���=��ʑ�c�O�����-hB���[���J���?�p�3}p�1W�~Y��-fj?FDT�
]��̖7Qª]:'�^��LVNf�K�!�øX���@��0c5=V�.IY��D�>��M[#����\�?/9����|+��l�9��s?��9ilP�˕�O�����1�z�s>L�dI�
�2'��P�����++O����C?6� �#��n��9)uT{+�R6�/�d�@T�����/ч�IP�ڱ�mD����H�N�Qfh�a��[��#�F�»:���)KzyU���}��6b�5�-���r�Վ� �'*%�j�+�ccx҇PbT���@+�9������?b?������Cu2���6c}�9�x� ^��.|��%� ���ANK��:��W���b��D�	͍�s��
�vL�����p<w:mP�����Ţ����빛����z�c_�\���z�f���Nfxe�~w��=іwO�0P)��4��;���4t�Rx�}�K%�2�S�l����o�:}&�Қ���VD�3pɤ	�1[}��r��Z��Qe�-�7&a0j�t���]
�g#Te�A�V5�
��,+�k_d�yAܠ���tF��/���TR}���,6gd�.�Կ';m�����C�K"�uB���%V�͐f����%"Q=6�V�k����R�}�q�r�N�+���y-Ld�,��#�@"2T]C�¹{���!��.���_���N���Ƀ�d
�=O� ������o��@�E2Od��n6��u�\�ཌ�!T��׹�7�Wk�׳DQy�!Ԑ�i�˽=�w���pz��f�3�)U�(���wC�|$����k���G�i(#���,�ʬB�W8�F��E+��/a_��E<�{���E�`�#�b����W�4<�P���O�\s���F�b��3�
I,�^7gZ�����nسX�zf��o �Vk�䢜*�S��	����=V�=���H�C����a?Q-T	�X�e�YP��.��6�,w'j!"�m��~(Vb&���j��V}�S��
k�� �9��Lfy��ڣ�D�s$�QD�c��OIS�t��@�A�=o]�&N�*h�5X�L��������7FG?(��n�,i=�u���{�a�/�$��Jc����w�b��T���x1��|4�ER�4?�U.E �Ӝn5�p�-�Hc�g��Q<a7��o��6j����
8�.�JW�����s���OPX�q�!��q�Q�J�/O�<����R��SL��sm�z��,]� =�$��U��-,uсQУ���	�^1PM��+�$wro���~���5�+�+��_
���:ٽD��P䋑 mx�#�O��g%o�cD0��ģۅ�R�Bm%��yI~��Xqby�����=x0|4�:���hi��$�Ab\5y0J��YV�4|�6��>gK�t�-�Q�?r����I���G��	D��u_����v�1�C%9Z�YV����#�19�W��):Bp��~/V�U�Ib4l���=��TyF����J7�;�w�]��pM���c}T:9m	�[���Ec?eŜa��י'0@k_��"�zz`�kn{t	�3�[�wIl�s�D��k��N�~0	��K;�� �s�W0�����Ŋ���n�֠-?�{��-�:U�2?��UT���&�Z;�8f ��p���	q�	��d0U�QVe���#Ђq�i��[4�-'tL@���z�}%-{��{�d$�fRn�.p���\^<ISLPU�*3j�rfKw8�Ѧ�Vt2x�c�K�M�+�RM/@��1~r�׆m�\kۧ+L�?3��b~9e���o"@z�#T��F"���T(
vY���_��B%C^��VW��u�:�(�e�����fV��n7�]2�۸�MqT;C
q�B���o���s���$��y���K��_aU7]��N �U �E�;�[�Z:�6���4���=��@^f}�s�W���r٨gJZ
�q�&��v>f�����s��Nv/���,�i&�%M,&�� RS��F���Kv��@d�?�'�G觔���X����`����K��#�Ҁ3z��%�ז=�.E}XU��:�	]�L@t����LЧ��Cok)p^�Z��\]/��p#��<�z�;��*�y%2R�5�ġ ���B�ٍM0���)Ϻ�:ӳ�x�9�7�27K����|� ��bCz˴lZV�Q�-�J�B���t�v5�6���#��G�l�T�*5��dq�o�F,���V|��
E��x*��㠿Ig��5�N��#�cV?�Y+�}BF�W̃�I��X^�(���U/����f�n�a[��4� p%N_�O����Ӫ1��&�صQ� M4����B��a)�D�R�t�B���"���i�h��ג3!Z�LU;ضk ۳a�)![�?��E=@�4�Y����/g%b}@e(Ed�|�c5?�/bs�~�s
bSA�-옌 q�|f	C)KkI���8{;w��pY\�=jISU譝c�P��!& ���eW��A��y���
(�;��S�Q��x[��Y9cz A`ZW�E<?���A�|��DC���+o��_{x*@YJx�2;���X�!������#x��P�}���H��XD���/=%0x�P����Sᅸi�T-���*I����h��@�T�$o\�֢JZ�$�ɽ�!��O��."w���w�+�O�|Ţ����x�vu<��֯�X[�AC�N#b$�
��5�m6b�>˷�{&��D�cN�� +��!�Q���7=���ب�2��r��',���>�x�^5lÎ�8�WQ�d� ]l#T�ƐU�+���D��en&�2�s�NŹ��ƞj�:�Ʒ�*X~�}f"�oӄ���Z8�9�x2ګC� �KS\6��{��&��DH�:��?�=0f�ce��ç8m���g�a�"�d�ĒZ�o������Ͻ�E�c����.�=������2[�G�e�l���va���4��%~�.��SKYCG�t5��O�1����ɟk�h��+�혅E���	l�T��H�T康/\珥���`J�����(��=�:�	��~���V�Z�x�=6�#V̵�7���V��r��S�x������f"�� K����CC��*lp��4�����R�H�4r�l�������C<:7(�	4p����pP1XA�X��>����z��A
UY���c� t����^T����F���Ө���H��c�m�ZN� jF�~���^�"F���ᗝW�ٱle"�� #s�"�6A>�۹�Q�uFV�=l7��n�Ӱ���z�`L�	�_��"���Nb ��0W
5�l��B���U�7�jWg��b�6PIT�Ok"����?!�.���2�{ x�#k���T
��r1"�݊��C�&�0�K��B���c>}Q�Z�Ņ���sI�BE�e���L�%ۗ �O5���`�O�6F֫c�+^+ʞ[o�{Q|Y��b����RY�^*���$�(������4����S�|o��v�r˽ g�:��{
u��!�C�𢠬�b��7Y�#cV�k���+)AF���V�{�Z�2���:-��RtE�KIU���wr��m\�u�!KU"�_B�"�3�dn�&Z$�
_�u����&^&��/�'!PVڂ��ļ�Z&?��%�:���(�(R����Wo7����	"�=�Y�VǠqL���m���&~��c��f��L�P�|z�f�N�������x�/����H��LC-�[�?B"Ж�'����!PИ�"��<���0j*���Nq���G+痉PڴQ����� ���x	+l�!�9��j�G��ل&�'-�8( Ϟ�&b-r���܀�6�S�5�ZK{�u"d��)@��*g�80��e���� ��[4���#������4rN��P���>D�9s v��x�,�^xTE�����v1U�m�L.ZڋK1�������;t�6�!�"ۇ͎~�Vb!:rfR�x�����	Yk\&���^����>Rvkp��}��u��A�U(�����}|��z�Z�y�H`j�Β�}�]�/C=`��Zc��/��x|��$y�|QۮzC�bӐ��iA�܂�)��4^�'��ΆљÁS�d�+HW�-[�XA�%S5�L��9��I����þ� ����Q�U&&��J7�ݸ�v~������B�$b��E�ώ�zg�)-��ٺ�!r�5�T�䌕��M�(��sN�;���"Ο��w���<71���1A���$�9�R���N%���w�M�RV�_��avX�ү�y͜8��ݎz�%%����&�c���@���v�"�M��
�!=�1��<���*\zi���L�*j�޸�!����9�*�.@�s��xr�~�ģ����G�ݿ�����Np>#�t4�oT�z�EzVE����������|*>ح&�����LQ�Q��.��Ϸ�녏���HF���f��ѡ�����ۑ�E�l��0l@"0��䵣�������x��k���x��O�?PC�Ps���4����9y�e3y�w!@!9Lp[���~�
.��]��=����H�jc���M�7�atS�il9|*"�^�]�/i(�,Yɐ�����`Q8�l��{����u����F���1��?��8��{4���d!�D��֝�?|18�G�sM��s3�:����PX�sN��R)8R�B]��1�{�ϛ8W��c�Қ~���,�jI�����P��;����%8�PzJ1�R�o���I���]��¦9|ȳ��"�;s4�πػ��8C�����o׀�L�zߥ��/���k��{E��ɺŁ�^C�H���y%[���J��e֭wR�����:��-z�����ny��~�sh�es�l|�}�Ɵ�U-�vME�����F���t\�,m�:��J�X]�Ļ�x�#4|��+>hˬ���\"��"��HTHf��I��flE��y�|��F�x\H�!#��i>�
?�&��p	Ъ�5�w]���c�*�] ��	�3�(�!K#��z����g��\��=�y�DM����Ryqc ������v���44H5�@D���?�΀�p.{c˾h�\yC���tBHA<�ꦝ�U��l�Q�p�#U��]�^��4A�����:��!U���a}s�{E��<'�j)�5)��]�OtQ�ʅ������vE��6;F-,辮�Vt|�)�*�bOM��g�{�F���o�p�ݺ�� ����H������jO�mP,^J������p�īcu O�'q�J���p��!
���	б�s�� 	���3H/_+�Sx���7D��b���� ,��"�O���@�/md�՛4�o�9�<p����Hg'��P>����&+��[�8(x��vy?�unv`��&��6�#�I�<�e����q`�D^���VJ{���V��dj\���tK��&<^U��d�c��:�U읣�@��!�Q[u��r�Ǻ�dn�����,w����8�$`6o�R@���bk]��/��>|�J�O��s�s�$;X4��m41dd�͸zӞ���U mpf�ȷ	n����p�ct�Z�ٜ���	��b�UAw�_-���%��^�+�-��HUzf;��Q�l�k��=�����b֦]7�c]=��C%��� �(p�%kIg��1 "�f@VZ]l�ǄV��{ɒA��Q�R�J��*���A���8����tY�:�s�W\p&׈B�T�j�o�F����2�Xx�g�rM�s���`*�f���C�]�]��*q�ĸD�@�������ZV[��ƛ=*��ƻ�z���#��0�A�R�	�����@�+���OF}��RH`�����&{(G���xK���U-���/��?P�ɠ�"ݳB�Z	��m��FO��W%L���3����Qj��M���_-�p�~��X0��	þ��۵�3<��H�3���};Þ���z.�Ķ�*�T�x�W%yB^�~�5�eP}����K݋?rO]&���xQxnvi�m�# w�Ɠ�NUu_쯓���x��Y��iF� W�g,:��V�x���."Ncy+�L���1@�@��}��}�Ε`��+栵1A���X���DG���K�����YM�;؄�bh�)��E�d�ǎ��	'���N|Nb��3�a��x�c2�,-b���sx��X��Ъ�%f����)�/s^����E�aW�ةv*<۝=��%�F�6M\����IW�Y�����XlxVHYEB    231a     6f0���Bc�A�%As��G����t1w/J ���y* �tTy�I>Mo�U[F��VQW/�bq����d0�	�ߝ��l����cwD���a��y6���8���!U�F�H z�f����+�ڟߚʽ���9++-/pZ�#9�_��Ta��۰���'�'W�6UkA�=v`1�J�f=0ﯙ���b$����ƥO���gw��$���5��P��g-�I��mq7����J�ޛ�O��ت+u��w�)��J	(1h�;e-��	�b��� �&�m�ܾ��R8c��I:Y��gЩO�zN�a-��1���mk|�&����;� /�L�w^��m
��M��Lt�	�v2���F¶K�������B3�Z��`��_��o�^M�+���ΜO }pP��h��Ǟ�ZT��"Mih+�n1A?�����*��F	x�zk�Y"�'K}��xW���#�G9��Si�4׽�_�yg����y�1���OH��Ur�+B����8�
�N�cl�~G�)���>"�稍�W�ܽ���r��inP&J/�D�*�b���Hm� ��{Y��>z��=��`2�ܘ��q��[������g��1�QY�I{���Q
H�/j5A��^[�4_��3l��D/��d�x7�s��èU���ϒ-��G'���[|�5xsZ�[�/��h(�`�+��)��h,+Nmg�fZ���ߝ�k���Ss��L{u��G/��18읦B���L	 ��S�.����m���I� ę�P+M_ϱw�#�&�`�����g��WU	"�i68��f%��Z0��{vd����Ț"���~�Bi�10<�9����S4p���0�E��ts�>	ts�rJ��K�^Z��Vh�#���QX��y7��ڔ��)�Id���	��S��T7�(����R$�8���rvO[!U��ۓ���n�N��,�d�2KJ#��5�߹;_�=җ�)�W�A퉼�����gF0|3f��VQ��L;a��>�o��C@L�*C��#�b{
��)����g��ݴ�����%ぐ�J���
63i�A'��"a�M�rJg��r)��mYY�^Hlmo���e/� ����a1[5�fU��$��ߴOo�;�V�J�9W%>���=ɴ-�\?!��,׵Fț28|֍��&[��݊�0p�r���T�I5���jΏ�WڛA�A�j��Qc�����Q�����2'�s�>2��]�����#*T�liz��\���^*~o�����%k5>p��8:F�YW��@`��O{K�pz�1^�{�x��|m�d�׌5��p䖓T�F}�x,�֬�e�l��2fK�4'�]G$�S���yҵ}h�'ݑ�-�����P�3:�����y;*��t�u�>����<#Ŭ�u㘔�Hv������}�o^vct*J��j�+sG��vu�縏r6B(�K�������ښ��R����Xg�'�e�.�Ɖ��z32ù�ԤÚ��񦾈^��(�c��SM48�R���j�>1�Ŷ�;R�1������,�+GO$���M�.2�K� \A�r̥��'?BW<��2e��f[����Hk8"�%�
�n�g�Y�JR,����jT.0>	� ���^������=B��i�f���^+*���қ�z�($;Ӳ�Pje��W��s�����NcF�v7��
�N�h�ZK�p�^�ۨ�u�E��A�D_o������n����*�.����� x?
�v�r��x����A��nYCۿ����);u��