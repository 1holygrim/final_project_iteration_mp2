XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���)zP����ҙ�j{��~�S�W�O�\~0����hUk
�n������Ġ�$�`�1v�H�Ɏg�T���`a)���1I�;��0;9�gN�'��ᇩ��=�)�Ъ�/��K.f���YhH�9E����=��	��f�As���Pv���nQ��Ӡ:�&! ��͡�c�� �P���(9�LDϗe��k��dA;d��`���o�lJu�CYG�V�LB����ᆗ��n�݇gn�g��o8�#.�dF	 z=��EG-ݵV����a	���){j����M�k[�N9�	�6q����]@�y�\�jlk��c(Y;w�]S�d�Um��b�T������6�q�a2��k�!�]�!2�,���1nJ-���<�{*���ޣy��LP>���<��]N��©1��.瑰�'u-R!��F�]��L���/��`�RZ�6�<�$ .���w���������Y*�jX�����ז,�m��xm� �7��Q����S��
����{�_8p�����H����������h	|��L��.�g���V���Ǘ����`�U!W 쭖�r�f*�w6E��t����M��u�
��C�`�K��H����A7��,o�|�y-�|���"��BX�~u��U"B����p�D�[�T�g�:��+�n]�}�c\��a�6����RR�W�c2	��m��]�)�r7���M��+� ckm�Ɲn�g����v� ����2�׳W}��Z�3@���
,�
ϩ��.�6�����'XlxVHYEB    fa00    2040t��B�&�@tyF��	�t�c7�����2�1ѓ�v�N{m�wW�	��L���of7���:uթ���L|2 �#KLt�5Hh��/�Ԡpp�ktJ ܇�
�h�2u�v���qh�e3�$��R4s�i�.�,\�j`��٥2�t�ip����W�Bp�0��V��Us$K�7|���K��Mu�yoaC>nT��Ѕo�U����XPY�����]+�P��{���S΃WI_бBYѐ��PhtI|�� ����+�aAT�
. �V�E�P�&�<݌��c���&{!��[���o*��C犘�8�:���5x�6� �+�u�ʛ��9ԃ��_ x�$i�7ˋ����2��6�N�8+쿍�~�4�����=��7W�Ê.�~�3\�>TZ�ex6�Ì���8[�'����]��yo����'խ�fjd�O<��������\|�VYWO�l}�j*H[���xe�%i��p�D�B���ƪ�d�3�YZ�т��>��ID�G��-/�����*ÈS�Q��P	�L0���1vE`�\�M�P��_�SLr([���)ص�va}E�N��m<��B���Z��d �e��A��y��S\f��}cc�9¨��?����v~BDj���M�b��5'���bI=`&�i<�m3Xp�[rR+�ɤ0U��J��!��G��	�������JR&���e$�7|��0�J4�{�1MK����e�8?4{�z����I�mҁ��_-���1�@�[}{àk���h6��dsaz��6,�9Uʝ�E=fBWJ<�V'��b�߱�O��8iW���`�:�-�jF�ܹxr�_,��U�	�/�����؇�Xv40<e�!�xY��T����^M�tm-H(�ܣ��սR�UnhD����@U`��r0�P�Ш�_Ӕ�RH4St�zl;%rp�~I�q�������b!^�>a-s���L[�醬�;,������d��I��q��L��?�S��}�Ŧ�d��歝9�q��3�`�ԋ3�v�8�=͸U���3�u���:�p@}_ϼ��;��7�&�|j�����O9��5_����Llol�]+fL��y���"��W��e�3����'9���Y���U�עڙ$�j�z���Fؓ���V�)������NR�oIg��3�C�|�gAF
�!�S�F�B��1ۤ[�8�D�����/Kw�2����-ڳ03#�&s�}�H��I�$fգ�)/����/�z��WxPl0�6in�5�펩_� >"t���TTd�x)�!��D��."�qR+�M��
P3س�Ѧ�
~�ۄb�Wt�)�Q�uN�i�"�V�H9꠭�����P[��o�����ga*e��p�JDl�@�Nya6��/`�K�`ŕ��O(��� T��]맂�n[��Y��lv�m�E�M *D��%�3=��d���Π���9to��+a ��.�ox6�\�уWr�F����?fm��&H^,��(ٟ����9 �ᬱiǾo'���?߲wj3Q`�Q�]�]Ӕ�)���)�W����(�W���c�$��3I5�5�������ͯ
d����g�[c�Be��-�V.d��$���/��l�H5?�qM�ɐjI�8������*�Gu�����L���!���tԗ��nzj��G�V����x)�[����QSn�9Ċxe(C�p�� ��w��S܊2��n�7��֧�6��(��k4+��E��XU��|WE�h�r�zP[s4��i�ƴ�(��&���~�WeUn��Bt1�y�m�%M�Х��)"��"�Ben+��L�N�e�: ��?��Ʀ�oإ���j��@	z�=+��}�P�F��y��s:��x8*�[��7$v�M��y:R����n�`!c@��D�~	��V�����*� �Q;��vѕ�e|,�*Y�%o�9B����d�0�Mk�8n6�0�-G ��n��#R�QI#h��s�f��_K��v�WQ����oE�7(�HO#��,���{i�Z0{�Ћ��U��:��ު���S�'q6J�d�� �(`He��Tgk����v��든�^��z�w�Rat�p��8p�������β��2��(��5�=��:5\1r%t�4hz�H�I���.7a_��7��Bp����x�"[�\�(WI���t{�g�����	�_��� Pv��_�]B���1�3����D"�S��8w��Xx��5���5����@��G�Br\�핑�Ǘtr�Pik{iQ���b�C{��z�i�,aj��}�iy�G����>��,���[t����������hU}6�m�����s�j�!Z&֠ϟt�6(�ⴀ��os!$�Tu�\rd�[�ǭS�k�}�?4�5�rC��[|������k��.UDĐ=�(�;$x� `�!>�:�U5�^H���{JNp��n�Y�<�w;%Z.�N1����ꦪ�l��:�_��d�{W.�4�I���l�с�\U=����깩p�۾�t���p7@��1{#ҩ~=�D���ݨ�Q|Dw����D9pI*q#���lH�ɠ����r��BO��]mGr&�|��Lp������aɰ
�S��H���,f��%Њ
q���"�VBvR|:=-���)���<�Po�x�
g���L��@^'��E&��A:�z�&k���R9"+��4c�.��!�v�R�+f����W���]V��RP�т�'I��=�g���w��oj9��4��,u�6��F(�Ǣ`X��T�G��D�?�d�D���lh]C�usQOg��z�O?�N~YWW�s��������i(��8�=��{��P���ˮ�XW����������<���ֽ�W%�hd���8k���6�p�e��/�a~N��􍵒24ϊ�l��`�e ����g(^	�ݒ
zpf
/�OϬK�����)	5�n�<�L �e��gn�-�`�GV;�Z�Ͱ�1�t�h�C�BA�$8?�����p�ߪ���jm��>Jo����0kV�֣���#C���}�(��D!��t�|�ͥ��	V����&�I���U8����[�c0�nWXkX�a���l�E����(9y�0�>��򑶁��{by)�cfσ�ق5d���E�a9�lL�$W��# \��%�j��oe�Y��J�'��ή��,o/
�=�l�^�7q?������!om��Y�󃴷+iGV����ċB5S�B8����L2$��p6k�r��aI2��pō����ќTkw�Vc�IYO�m����ܑзc�\�+Q��twE�e��|�!��*|^�u����XR�Ɩ,*TN�ͅ!��PS�Cۧ[�aAyA�h^�T��|V�,y�Å���+B�c�pn�i?mD�I	,�z9;�7�?K�e�$���q6
������hB�,P�t%a���o�q��S�.!08E>֭ �{���U�_@t(8��_�i�j�4�L�$�Nʨj��I+t�ro�#��,?G-������!�p�]��Y$�"�M% F�hb>Fp�~���,d��w���׭�ү�?K�HW�G�Q~9��;�?�&/5�P�,��s,�2U[ �>���������5� )�"9He�;#Hg�p�Ag�p���s�D}K�[b�y�<�B�e9a���T�5�Cm #0����20Z��胑�"��E�S�Z6O�6��˃ &a7�B
}��h�����-��>������Pp��k�g	�J寣8Uh��$h�,S?��]�:?:��;������t�Gc
k�Vt�w�Ok�Yq����y����W�G���Btl�����v��u���d���^�Zm��H�{���XB+�m���ꕟ;s��s�$��ooĨ��}�f�g����t�2�vMH&�w�f�MfŦ��X�s�5���:�����aD34d�vK'"��v��$ۅ�g:\�(����L^�L��Һ�vh��U�!��e�a ow�P*����o�	5��m��	���	B����O})��%u*���hR�Y�0�^22�����ͤNs�Z�a��\��`����-|�V�9��L �����R�1m�>��Ε�`��%�ă�0�mSy��7C���]�;����/�I6�P��[�w�e�Dc���3��T�5۴S}���	T���Ƌ]9B@�e�,ۋlP�n���̎��o����6�꬐��z\�#�KU��F�ec���&��u�O;ܼ���GX�L�,��(ʈL�;���͔�zՅ������F	��x��m���P!T``
k~I�]IOzjC��zG�]?}�F��\F/ung��8�X��I�gd]l#x@ze&^~F����tW9�͝ PB��=qe�r�_y �a##^��ٲ��+���������t����:+2�*q�-s5(d����+V�� �IPab��"���7/��pP��m�f�|�>Կ��>>HDA�l�Q�*P5�c���Ԕ3{3L�� �DMȪg/>۴l�A��2@@d~Xs��a�&�m�۸a�b��&u\�I�f� ��]��\*!&}��Ts{��4�dp��[c'��D��c�#��ɻ��s`�*E�g�3�\���:�,%S2	Jf_��7ήwK��f��m�]�0���ӛ�l7I���\���06���P� ���4J��5:B�/e�	tZ�hq���w.x�P}wb���������ڄ����@� w��۞7����
A��迭�ҷ7�s_�/��!�+H�x܈Bx��x�-1Y�>W��^S�n���kϿ�ĝ��� ����Q���Ô���m��!8N*��ELj�1#u�(n�9��}T�i�����b�w�tl�{m���B}�a�/�eK}�*1r�u�o�7��8;���I�Eߞ)*fl�,�8�>V�O������}>�7<���^�������S�4И��4虣����R�c2��pJ�����:��}�
qG�e%J������p�"��k~�+d?��ftB�{ J�-���w�ÎW�I�;t�D@�������(P>F%=*Ǝ�p�*\A>�gd�T)��b�f����&9<<������vO�o�t�<ì3.!lI3l�n�;C�_��J�y�y �+�	���w���Dl��K��@�9����I�+5rW!Ii��x�e���Ct�L[�9�h��2D�ˬ�Ȩ�ti�O/��h�F@���$����&4/�x�0�) 2�
�	X���D��,�K~�d\�'GM �a�/3y�	a��Sqn�<�]�-"d�yc	�
��V�Q�� ���Oֳ��l��T>*ʞ���Lx������簼e
cE�v�K�Y��]�	�2��!T�u�Aی�8	��N�=�z}?�U�"��0H�H<�kf�≿0�ͺ�k/��K����-ʊ\��
�zL�������Iw3�K�H��Aq��KDӧ�@�\<�D4��X7>j�� �kӲH�>�
��E���C�vU��A0 �;`��bQ�g��-���1=ߥ�6ƭV�iW���t��;8c�?���fw)2�oi�B�YP1�_l��:�nm��y���� ho�;���4��&����b6%�W^
FwW�n��U^^)yx��k��I٢��֤e����������p��ɑ�{z��u��Ix���4/P�v�3��e�b�uX|,�8#x��8����Y
���d�M�٠\���|��Ƥ8H](t�K?9E9{����u��e�C���ɘk��ch+�ͭ���[���+�3�æ=��T�����x��6ď�0T��@=[��?�T�Z9G%�>C�1�!*��'���"�ŧ�A���?��ox�;,���4��JE0����5%�����R�CwF��i
�懧�O��R������:��Ď(� �ˋ�#${�S��o�}-��F���RS5��`U��1g�ע2M���ճ�H�����$J�V2K��̽)�9!��]�^�����W��Al���X����>N??z������m��������D�ش��+�jH�R]6zV�/��.����6�X"���%6��[ʤ1x�x�B���0͘��sk$N��)/�i�ˉN���+���KKЖf�m�6�-Td�/]<�����<`+�~.{��z��Ee:L�"D�#.ݦ�뺷⺄����3O�[�I韀?���R
C��|��4u��D�-G���N�=�ьb�������i8���_y�y�����E;�$��{���Jx˒"�v�Ĥ.�0K�Ti�є�.���nܷ�ə�L�n�@��/8$�ok1���q�oXl!�)`l��cK�n��5J�]��~[q�]$[b!��VԷ���6*�F�/N'6RX�'��`0Y8��WVP���W-��wlM����3��R>��8Q3e^��#eg�}<q�>���߀�>⤅h�?�ip}��	~�0�X��c�!����[7�J(/8�Kup��5�#�<Z
�<��^��v^��Ů �-���4wdt{��1��:-����ü�x:<�vV�
/���7S�Zo �s��!v�y���s]Vêo^Ι=�>���N�D��s�3'<�U_aK�4:a=�m�h��V�߷�n{]x�=����������M�]d���S�V�t���Dh��~9H"��3�w@R�*�3��ML�U��@D�~n);��nf�+��������\�%8t&������!�CU�C;Y����!� l�Tm�n�Om�V75a�}��e�,v�h��i��:Pf`<�iK�_�"����Gq�R��n�VRI��`�P�~{�tg����,ǖy@7j��%��ܴ�l�$�n��T�2k�����k
&���Y w5�.� �| #��O�8v�[>;d.gL�Pt<������􇴗���q��,��Q���������{�#��
�g��L��a�8�0�Z-L �t^��I܂�����z�)�m_�I�XC�Z��Վ�=�$�}I��¡�Z�/���0_���%��c�\��w�� ���({ۡ�8���B��p�=˛М��ej0�N�/>]g�Δ��E���CU�ݡ�r���o�e���K����hV��e��`�R*���d/�zkZ�u�ȿ��;�m7�U�$�P��-=�W�޸F�8˭�u�DxE{�4��)Z�G��� _X�q���+��6�R��f��m|�?���Ư�@I��dko�c\˕�UM��S
�kJc�a`֖a��6��iBH��򢂜ج9���S��z��r8��g��bF�mlyNhSP,��3���a���y���ĩ;76�iX^2V+��A����� n��ZF8��i����;����U�۱G��1+v#��[v:�}��%o���sn��K� ���V-�g��M�6{���Xw�;ҡ/��p	�3�Q��e
�х�����ǰGZ��c�k:w� 6.�È4�|�h�;��j���Q,^'���ļ=G���Nq�b���B�ނ�D�KҞWL�^�\�^��Ж��IuY��+�E�>�}(4�?�¸ڧ��v���*'�~�q@	��	>癥a��>LkI��'������f-�����'��9x�SQћY�,� ��F��nM��]D������:j���������?�f?]�ھC��$K���Y-�ң�4n��4��h�b�q�(�\
�I�8��9P+���n(���+���A�+�^}g����� �ĘN]����9���b�7�ܵ�F�A+w��0��
����l�!����@TEm��݉��AR�фNmh��pX��Q����q���[���5AxP�cNx�ް՜��T�e�J�ss�����&P$A�bB`:����1�[Z���]͎Ιd{��%Y"�2>����Sh����\���<�}0�"^B�Q*�lv��$���
� c��{}���0Y��y����c,j�Q�or!��ypC�e��$�t锄{8~�x:���[ZJх��ً��dϷ6�G�%5ڨ�!/��*����QN��˙9_�Œ��5���ǜ`D)oVWO�h��ȺF���]e�M�;�P&\XlxVHYEB    4f62     b50��բ����$����_�xNV�k�d���o>gG=��J~�Dr����ۨȪ#�@e5ı�.��t+���1@N8uZmb�(q]�x��0�yb\�� �a1��5�I��+��dLsچ�v�=�C�>�;����@-k�/���+|�H{ubw@�
6�9�1l�	��03��P�1`��AL�����5��������!$��\+�j!m����`~t��0 �H���2����z<x7����xJ�������)����ˈ��J��gG��}�nL�+C;���k�\N�n�J�`�������Ø�����b^�H��I�T� �����*�l���g�ѓA������q��w5`UV�؄�od��#�����k��Gg��Xvs:#�������6��p^�9�/6k�b��XwI�x<���+s�U��z���y�F�[�G��
�{���RA]M��k���}):��{f��+�����8���I7��3�Ԕ��އH�(�Od�k����`�y��g�|т�o�zN3{�l�F$��.���=��R�.���>n��)g�ƨ�r=@��u~sk0�`�9�:�8�4	��Dh�&?]@H�]T�`V��锾R\V��{���C�uy|ip@���Axg�����V�Ǻ�E���0��lℽG^�3�o=^	/����8��{�y���[p��Q�񇾹�R���T8�l��^�^G������6:0��#iׅ�9'�H�& |�/��|C[<�=�>*>x'c�Ʋ�d�*ڑ�O��������n6i��]���ϫ.�;�=�/X��^B��v�2��=cx���s�&��Y���D�Tx�l��[K�
p(z����m	-7'�R:9#۬e9��\�خ�dv�D�/	P8�k.z��BK9W�����#/�c�EM5���7ɐ�ľ�XN��@:
�XF�5���׃��HqZ��E �~� "�TKG	���K!��,�%D[J�#�%��������sM9����s����}��c�f��\[���[t�.%�~"��v�=;NU8���B�F �<�&����|��r�Z%�-�	H�9�lH0sF��ܩ�׺R;8\Ӯ�$X��4��D��m��P���Qw����R6?�g�����A؎���W9����GI����- [J��X��+�p�m��8�-�!	������(i��Ve�('��DcY�ڐ�O�II�3;4Ey&,f����q.^��n���H|�(Z��ʳ3��X��㬦g������O$P��(�mFYQ�D�_�Ŝ�_�P��t-�f�Ų;!��T-:�Qa�	Mm��2�>rr��S1�}tG�<[=��:�]u(Ə5������K�B�pp�g������hS�t��XO,��F�}�p�=T0�O3�3���o*�K@y�@"BQ1��u@�^%�� M�/�Ʉ�%0���{\zR�F��d-(��WE�mY�:K��bѡ��^wK�.�L͉Ig�rL���&@�=�M�N�#Z����7ο4��K\.n����P�ws���+�&�Hh�����Nir��J|8#$�;��ym�8���"�k[�T�ΩO1��K�N�Ʒ�ݑ�L�k���k����0M��� �?����pq/T����9�}���_&$�qe���#�]����&4�_7�F�����udo	��t�:0E��~�C��.�
�Q�H�8�� �(s.C�*�­eR��շ�Ze��M*�Z֜�r��6ɰ@��^�^ $Kc��ż������^'`�-�Q����M��mz6Ҷ[�wl� �JhV��k� ��]���a&V�V)���ɮ�)���*�O?���vj��V�#�h/�;?U�Q�-�UV�y�'�ϴC!X�#�1��y����1r�Wm�$C�m�3��&8R�P��%�(Y���J����kA�P��Oٞ/vl�';S��h�
�S�;ޒ_������pqV��R�O���F���DՅ����z�&�/�<%MYF~��Կ��:�s�����4K�I�#�?O`���NR�t��x��ֻJۡ�BY3�'ؕm���'Q74�N.�2��V'Su
��A��1r��	�k<�#\냯EHt�������Ѫ���"}������(s��@{�:~��?
������̞� �� �IU�-kM:@Ț��B��P��ݙ	������N6+Q��VjY,���U,k���G��{�4�Q���{�.�W.G r�4Ba�D�1�z�C�Ux�I��I:�fI�����\���`��e�z^N�����H���ꑨ,�v��=����� �(%Wh&l
SY�-��{B����a�P&{��Q�6�I��R��e:�X133�+(�)�B�2ts1�:��n�/$����Q���jc\ �ޏ)OA-�-]�!W+��MI
��U��k���O��<X��Db�p�lB����>E<b0l|S�oM]��flk5���=r�֐��#K<+E@�j�3�ʱ�B�l���_fwSJ!����z�4[}�K���Um��T���8`��zD�kָ�o�x�935>�'IhnW�0�;;��g�K$܊/�bl>�ʙ9��>��<[�3aR6�h�ͤ.��Զ:����0k��-��r��YA��nf�^��B���_�P0J�'�c�l��Wȣ}�k�%8��)k�u�at9�%ȭ9�� f��c芿�(�D���?��8	x�=��1����fL͏ǫ���y0z"���M�e�l\�V�������W���C-�^�T�Y���m�(��j%�ޑ�s��,�WDώ9�R�Y