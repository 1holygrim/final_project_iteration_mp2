XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q-;"��W��N��p6?}�F��)F��Խ>���R�F�-+��-k��L�?�F��
�ҵ�qF���
1��t�j������֭�ys�EmN��������b�'H)�LɔXo=���8�>ݖ�tBX��_��>��"��'�=���%i�ku�����[`2��1x%��w�ɶi�V�[=�{Xs��~��P+2�Y�@g��B�ϻ�5��K�ݢ 󤄪�jW������B��v�|p@��᪾'�Z�\�.b�����"uD�f�Ԋ�nȭ�`C�yڮ��d�Az�]�����k��L<�U�s奻ɈrF �Pǽ���Ú���սt��+�<*�S�P�s崍6'�20U����&��l��؊����1삷>�3��أO#�%IȄ�z�h&����W���Y���e�^N!�;_�j���oXɫF������d��تw >f6���pQZU�w~�>�� ��{���C��k�,?�[�����;�o=��Z)s]�}:��<1�,������!g�Q>=����E�0Eݔ����y������=B��컀A��1�`ȳ��=B�
��k[�]5t���H����8��#L�=�8�|*U�ie�w�j�SZ�qq.��l��w�ۤ�-{�H�^�xP����;��,[�]ڝ��QmV1��M�Ց��q�6^��u�LӜ̽�颜S�b���R3��H�����q��X'`�9�#�b��nM�� RXlxVHYEB    c05a    1dc0"�ܵ�;�Wɯ���<�g��iɹ�<��E��t�5%��)�7���� �H�<jt�ɯ�T���.�٬uR!i�s��W_�|;Q.��PPǾ�X�����}ah����V��-xJV��d�k�Y|F���vN��K�"o��]"�`��ʠ�;�a��К�v��{�k�y�!�R�umL�"�98E_n��@![�ܢ�:Pq�W�Z]�j�i��Ӗ@��	&5�޼�\.�~������|�����lʂp�:l��V/�Ξ��,H��~���lgi�s|�O���@��
�Jb<���������Z�s�k(w$�a���6�8=�	���Bu:~�S��;E��v�}� ���"[��13ɬXl�Ƽ�C �cB��L��9���8S� *z2R؋+���,�a�B@���j����+>��_��?��S�\�Td��o��z�E؈�m�W�:�h��dj���XN���L���ig=]" f�#ʼ�?4�_���޳j�Ld;�|�R5@06Z�p?��|t���T�r^����PM)]�@XC���+��#"kw�����ݸ�t�wy�V��&��Iˀi�ߎ��L�e7�?�jkZ��8'_���I�@��̍ϼ����X���*;�l����tC�ML�!<7a-��5:O��Un� �N0	
C��5���n���ߤ�!y#/~z�`6g?����8w�'�\�@��\��P���g�z���IQA��Ĭ��V�]nզ'C�i� �}��Y��s�;3B~�c�G~�BG���*1�Vuq��t���Y�w�|�����J�oE(�9X��'���[e�{�l��M_1�ytW�R��Qj��f!ҹ���v�%:��l��d��e���D9/N3J���|������3��w�E�o#����|.~z3�����l�a6q�~�c�h�k�%.}G9���g5?<��8m�0��v\�>�m�K#��'U#���h�&���!�	�� WH%��wI��NIŚ�N����Uh/�q(L�ج��X��@��GB#��oL!x������;�%�Q9�߼�������~����ī�t�j;G��"2;Z�|MHi-���Puf}Fm�G��c��e�o��(8r�K��O�2��}��0��	��|���fT�dQgS0�%Q�C�P%�ϼ��o%�| �tD���8s�����i�`Z�&E�+���nG���ʩ��P�W���B��q �G���*��Q#��P�M.]?R҈)y��YLP� s�?�H��}cP�u�յ�E��3򯰯|��Z��ݟ������	8�߇,�:�b��6�8��YE�J��H���[�U�9��
-�?،nm�+zf�T��7I�SU�A-��8�C�y�Δ�7��>mR�M@aU��u�e ��"̓��G_IQ�MWG��!�`��=dxbƞ=��#�bEǙ��7����4Lѝ[��#\l���w�"�1�ڲ�%����[�R����3>\Qd~3��v��<�j�J�\q��D��(B��G��<�~ L̾E��E��)����X�Or�;у��O�9��r�O&�!���=�n�e�����j$	؁�����?V�?W/�B�e����&��u�����V$�v	uȗ��vt6��b,y��`Խw�!�a%�f�Xe��ӝR֩�۝��X��Z����:�'^�d~���&k%�zK�i� ó*�?�(�m$N1����Do�o�)$�1�]aIbl;;$��L�9J���9���ҷxe�����G �1�3��E�Ϡ�wYQ���s���+<	�3���C�+��m^Ԙ�o�gZ�7	s�(W��]}4��DSl�!eM	��1�ʁfD���w�`������!���`��>Qy��p��{nz��->L��6�,�PcN��4i�|�p5	ڝ����J�T��Z_��>����r|u��`\��[K�l� p ��;�x��ڏ�YRB�X:���(��`�.��#�b����C�6e�ȳ2���>a����R0R/c`mBya�p��h�Hm`���.m͵c��;�E_8��sI�����`E��Xo�Km�e�N)��b��ȼ��R�٧�)��e��;2�D���8�sw���dU{�ZL-q�ub�H+p�x�/����9�gk��/VM��S�Z��C��^���WէG�L����w��L_P�W�-D`���xL0�+&��r��NPcS �˅O�����	��h) �g�gN�iQ$X|�Ƌ
�]���S�2޿����R�[WIH�L5m�W�_j\O�����j�f�m���h]K�/ms[Q|���✺�9y��uT����s�;����4���n�j,��7Ȣӝ,%Zܛ)�O�-�%��V�/a�#QF��U7wd�Hܛ>��y��O	�ٞ�3p��Έo�ċ���F�E�8��_����:�0�j��	�=�]j�#���(�U��j'o+��R�{y�)pڅ�H�_��dZ�S�QQ��A����C�	Su[ѧ��;�'��I��936Vǔ���a&��E�B�����
^�t���*��zF�j�so���"�fDF�2�����������D]�ԓ�Bu��=*]�L�����(iP�α�����:b��>��(UL��j^Е�����l�|�v��i݃�+"	_:�� h6��Ƽ��>r[��W,��qQ���cG]�j��T��Ͳ���-�g�#�X�fG���9��×�1�Ñ�㙝�yQ _�HKOg">���#���P�~h�s���)���=P�e{�����Q6b��p�"?r���M�b�����~�f��F�-3?g��e�Xq�|����]����T
�蛢����)��)y����B
^w��}pY�i�u�鷺1�Fu���q��	��T!�/L����Kv_�?��yh��Q*L?e�����l8�oCl��FmC^��F'��X+my�@�a�
���dF��Ɣ�60��ԏ�,/�Z�z�{ͫ܉��˙�+2�ǎ�U����Ӡ^�ͻ�S��_>F�6��f�pd��ΒbNǼ�L鉰ז.�/��U;�ȹI-�62�+J��i�g]r>�;��PO�=e�H�<��x;[�䚓;�5�`��~�g��e�)�ޙB\��K-ӥ��r�G�L���D��"��P�A� _+Lm���b�i�.���<�慰����П�/������Hh&��3n�^����c�����M�|�^%i��ra�(�B�p_7�<�sD{7)�N����w`��.�GZsz��/��,��l�<��(`e<�|R�D��陔����,R*��Bh�y���G��M���(ϊ�ԟl[�B�s��D]<��	�$?�$'XR%�P<��$�i�-��}T� �ϕT����-�e�S��)(��@S�Ec���M�4!��&���XHе��/'��ɵ���K��-FkɈ�G�?^�$�z:n_��>����o@�*��ġH,�G��m��*
A,����:���h:/�L�G�:���G�R�i,w֙���b���� {ϵ��叼l�S�]ĩ���^d��sҫ�V�|�Е�	�0���ƹ7n4��8a���d�aL���x�g���wf6�Q��MjR��i���H���@�׵%C�[02V��V��`�{�zL�_�E$n��˼�>ݙ�?��}��ƴ�gT�LXU�E�al|Z�N�ܢ�9I>x�&{M��&�D�u�����$>G��D�j��|�����]�r�(���Y��@��--8�E�mH���}*��:����Q�z�>��<���y?
s�c��y��&�M�U�e�Jv�~�#�N.�3N�6.�e�P�X]H�s�h�pE�:t53�+(���c�,-�;��Ӈ�ڐ���.%���g�6����>�o`�>�� ם���;�t�z`/�5��@�d� �*M��l�W�c��{�xF�Ll�p��©W�y�/���,��m�'P2a�]H�ux�Y�ݩ�!z�	�[���ݲ��g��-��*�g�����|e�l{�l��Q�Ʋn͍��9�zV��F��s��z>�Vŀ'����+I[��ˇl�O#%B�~m7*�3| ��bHG���v���C�yA=��C�`���U�<;^�5� ������s &XC�ym/9A���	�v`K[�����fڃ=�*`�i����1y{L�4v-$Q؀�N�,jg+Ϧ`_g���3v
4��ݧi��I�:�؞u�
ސ��:�� �֒�{0J'�,�D궀��=���l�ZE(?ހg׫;�Ÿ)y�~��D�bz�8���2���5Էf���G&�S�2�Ȕ����i���ϓL��D7�ކ����4*@S<;�i��5�sY<����ٯ��#��`��
�p����T��kgP�di�rU��uSٛ���>C��x|!9�Շױ�M�AH:��R�*���RY�.��4,b����� H'$��V����_�ah�l��@&� �'}��TK^$���SH�jn��'��YX�E8͍��^����d*)��vf��ζ*��fH��%4[��9E"� "rY%����JZJU�D��"��T�\H�B��Q���R#�:*��K�7�0$��' �܌f�Qe>��9�3M~|]�$QfU���2՟����$)��[9�ޔ,��7\�Rxϡm abU<��ǳ;����dJ�|B��\F��F֦e���Q2Q�|0U�H���Z�M�ǃ��J#ؽ-Ҵ��pܝ�@���`�(����-���à,�j�_�ξ�)V�x����kBH�g�����7��8V�W�46C�N#RJLn���C�\,��X��������q��T���:�ʳ0L���'<(	G3����>^!|�)��8y
!�ɸ&�!� ��7�s#�l����O�� ��&�C��3C3�7��9�?]�;/���s�����"X��F���g��G�1X���C�����ׁ_���-ᖲmfL�ˮ�}UĹg5ֈ�g�E�5�/w*8l7'c*�o���ʳ��v�U���X�:��tӞ5���s�o���k�,P�S:#�t��\�=Љ�M�DE�_���_.��F�K�d�#��8D�	x�7��o�F��yv���S.m��Dt:�b�]�X� �F�i�!a�W��!V[�8�?o��=����+�D�fq"ShJ:-.L����}���Hm�R�gX�@��<���{��z-�
q���`���*�g�5�N]��A&X�f$�!��1�1��e0w�������^�D�#�	���M�?�]�V�����x�]*C~�A��*�Ȱ�Ъ�)�9�W���&f��{l�i����hOv�/�=���*	;v�O/L�.��F��V��r0���hIOh	1 a�8�H���S�{8&sA�賄�����/l���-t�sQ�I�V	V�-հ�3)f��s2 9�͍i��<���5V�<���z����H���)	��'d�wuvg���r��P��(��\���	2�9���U������Wg��xC�H��h���P��p�:JJG��İ�C��T�Vx
p3})k��R_�6�7wr1̥%TS9���8�b������o���QK�v�m�k�Bh&��=�E����H�Ⅵ{�
6�W[�}-'	;p�Z�jه��Q�  h4��+×����A/�e{�r�t{���@���Ԉ����x{ű��Cy�BW�K���������!�G,��A���׳����\2��|#�1H#}�z�T��"8*{k�:�Zsiۥ��q���&=�X �R9Tt���
���,�ZY�u/Ngu�HgH��|��x@��p���!X~�>���ϘfNr���!��s���	��@(����U�A�n��Tݪ��J�i~�-�aK$OL���T0�[�Q��R���Ţ���I��>�����[�?.��c�~���Ű�"��5A��-�;"��M��.�@i�q��V.99�f�uz�t٬7O90g ��#�}+~�x�j}vk�&h����8T��;�Ջa��m8�&�o��Y�@'��w\Ts�yq?E�qRl��*T���B�eLA;k�Y��u�2Ƞ�a�n���_剳g�����V��7qI�쇥,���D�tb���K�S?ͭ�F-���܈�N���Ap��Ϯ��vR_|/lO���k�Ԑ�ߩ|�{擕���B�{܂���a��D�0�x6�w�a~S[���񤑢IɶY��pO�>>Y̽�����.�Oѕ�H�]�RX���R5�y�(��tDX����D#�c���P	ߊMK�\Ha�S*�90J�x)�@���ܥ3\C�4�O��Vp-��P����F1� �	X�k��T�r���pP���)��ĕ���tE�\�kX�&�y��rk�AW|�5�m�b0^_�,��Jwm+h�$����ê��ܠP��dp۬# �T�r��+�N��iIq�e2Ӵl�<�&z��[�~m�`g��H-vK��l[:[��q�n�W-~�&�(j�w����D�驧�VeC;�h�\eo���J�#��T@�肷ܫ��?�v��5-���b�aoZ�����eT{�J�|�,��~��bܙ<he-&(C�pa�xjX�Q�zMN&-���+�繩�Ph)[�b��/�92��y\��uk&+�:	�:QR�ϴ��1-�����?��s��
k^u/��
T^�t6� U��d!'����c)3fY��ћa:�L�q�t%��ʒ~��dý�������g��BӮ,���Wk0ay-�vp���p�8����Md^�`����y$6���_I�ޫ���K���R�)n���C����23F?�yR$n'���3�= #��Xd�!ީ	Tf�>�?�
t˻�����!�� �^�Tד-�j`�@��I_LaV�l�ӯ3*c=�4�q.�:Ƣ_t�8�ۦ�"g�75bF}��(qQ&��� $N'ڑb��*�1�o�c���!�47�R�:��O��p�X@������0R:�W"3ﲖ8@S�zO���,�UT⒎~��7�N�ކx�T���A����M�L~s�V��#*�g�d�]�K,�k�%���D�ta��#�+��CXc�W�cb��,�1���+lB�Ӷ=��W3�v���t�K�M� �B�������j��қ�U�h� y���ڕ��)ej��vz�����ǻ+��G2.�&����Ӑ�bvȎmI�{g��&��7��uN�Q[����ɹ�Y�Ae��ҡ1��|����2�ݰm���:�Y:���p�Tʧp���pI���G���7?g��)ozj�D�����OX���Xe�?s?��4���N]���ƃψ0;{���h�\�D4�;�Lq�q����5\�K\��6�e ��qJ�!���i<���*{�c4�@���֑_eR��Q�i���&��I`�Tj'e,��ovY$��-��9�9 3����v�»� L����F�cn�L�6�.�C�.tu�����	P-�)�jU�C>0��7	�