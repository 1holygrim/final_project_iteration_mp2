XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H�K0*�9��3��ҿ���0�J)�[m��:ia�q�M���}�bO�*
+F�u�8"�/w&�.~�+�����p!2'�H��m�,��ЃK�^}3�[kީ�1�#�kG��mz`S�_�ֿ�b��c�.��m����Mm�Ưu=���k�KL�qB�S0Xe����1�y��Ƚ�H����b�L�U6�1|���"��*v���@�W1�06Jqֵ���(U�6�7�'�E��u\�
c���M�4@Ո����U�c��Y4%�k�.�i �|�Bq#���#�:��O��(1ZBуxA�;݂�C���.�닻?]ri���Ք/֪��,|���%PO$҃��o��̅ �e>��GU�c���^�$��Eޥ��ff�tU����ۀ~�H����x0[�|�A/�bw���/A�B1��2�%���(Zo�_��T`y�u�,�$��$���X��K�
 ����O��,H=v��*�u@jH��X���4����n��V�E�)�H ��e���Hi�Q�ˀ'W&Z�մHJ���໭"aѹX����W�I�I�Չ��*z+�gT���۹� �Z��T�q%����]q�B���)]��N��iǩ��nSk��DOnS�Q�|��X�n�2Դ���z���B0E�k��M�߁]��,'{���;3�"���$ik+CxK����ۢ�D���8?���������%%�	vHF�!�2�r���NN�D��L������)�o�%SRt�Q_ʕ5�^���4����������yZ��XlxVHYEB     e07     680 `���H�(�	̵���,���ܭ&����z�c��#��Xv�¾�o�����gp7�����eu�r�f��ϳt��2��x���rk�e�,�D
��Y�*�(o�=��FAڐ����2p���9Y�ݞ���w=����[��	|xѩ�<�싀JM����nV��o �3�H
h����'��6�sa$�5h �( J���v�ܳ[a�v� �:��:4=_n��3I�k�E��`t�����ɣc��u	h�".kwh��nvG�7�<����j/6X(-�Mc�����<m���{<f7D�*
_SҔ}=�Q���[Sr�_Z����b��L�^G�P�r^wl^&:&�R��j��Hľ�N��q���lZ@�J�m�9!���a�,���-�UC@`��&r�1U�FB�T��M�����ZMa[dCB72��~����GVPC�?�*L�)��躞��ԡaQ~O]Rsj��z�(Vh��{bBA^ҝ��p36�O�.o'4��֜a�M��D�)����sXw#���\dG����i$��x�~쳩~�c�g�6�<��g�U b�t��YaSӓj��n��2&�P6�{��i�%������;뾻�p�k^fF�Ώ:�h���P�^di��҄t��~�9�ծ��e�2���;)�NWs�FxD��m!77I@ܽ�N�"A���U���B.��b���hiS#�.f������1��rX'�G�<�ԙ?��'�:_�}$���E���w��#}���m�w׶v?�.6gɨ�sMF�������n�����p`����:��:��⇃DDj���U �A�m�2C��F@ܢi��k�nWo�\����d�����{�����L�젯����Z�,Bf�p��\�-���	�܄]��.�J7��&���
�JE�MPx`���d��#y�s���9!V4n���T�uU����+sR�5N�1$�[j�>�D����OVt[*z mH6��K��yC��l�%�`�_���{��T�o���9�df�G;P�l����sX�'�8������j�+n�9�0��%pG����D�V/I�Fjq�^�Q���g�=����$6C�h)������}��j�]e�6��+!��ngW03�Aט�H�[�9)�(�L�"��p�=�����|*���Z���z�S��ّ&t�G
'�ﱫZ���T1��N��pذ�x�	3]ja�]�G��kJ[*��Y^��\��@tX"[�c-P���[�YR�BcG�8�1l�	�J56���yϴ�j�����N�����[n�
2)�E��o�
�ã���?��������)�eArw�O�菺'%�C���T�i����P�� /0Ml �����e���?�Bݏ=��ZGI%�^3�b>(�U"S�����;tpK�],N��Ob6�~%I�e�Q�Q�uk
� *�6w ��Gd'P�hg� ����k&x�T6�[�~�z��Kԥ�[3���M��yO˕�)r��G�&�dWc�>���������+S���<v<3�
GI�6]Em�9�J�`	��0o����z��4��	�*�Zr�����%�p�5�����t'�