XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���>wQ�=J�{��J�u�=g6��͸�t�<��(��	7gm��/��o=#-;�;�L�hl����f���7��v�1~!^:���m���&�e��G�M�E$�u��?�[�s~�
E
BE�|���Mf���j|˲�@s�;�B�k��ky(	S
"�:�,�l2{�嶹�"��������������腇���I(uYhǶ+D����L_�fT���k�kbí��fN`Sd�W�W� �&Q�Dw�@^R�S��f�lB�)h�˗p�]����� gB�H�ǖV�fb��ݿ��o�,���Þ�w�9��M�%�$���C1�G�#�man��������uv51R~��x�;��Ř\������"k
މ�Y���l�D#bG��b��q��X�O�Qey��/k�^�IH������I��v�@�U[<��(*V�3�Ǧ#%0�l�]=�R�;� m_�dw�2{~B/�N�1�ڍg����\�o^L���=��e�)��J1�^�i	�������4A@���`e9�i���/�ׄ��ւ�O.=��u�%�L+xʒ�|�ri�M��u������1��m�~���'���0j[�n�Û��9��`(�­f�qq!�#�K���B��8����v�B��:���!l'�p�a���O�G����P�Po��)�w��B
X��E��M#V$����	��������${dQ����D9W�����p]>��{�k{0�M�cp���XlxVHYEB    4284    1110��6��[N�q��Һv�<t�2��ou1�n�̛Ua�R�
j��a�b[��Lf���I�����������U<ı��W��1h��Y9�e5T�>��S-����?N�V�׾w*o�wd�����Q��[ɟ�\Cr�8�����y�0�>Ao��*\���4��j�2����Ɣ�_����K�6��Z�j|�$�5���?�l$x�/����jW�S�?W�ν�)�@CVi�c6��J�_��O�$����z�D��˖W�J̤�J�UYMR����uۼ.(i�d�w�r�V��8��i^�mC.EoUOH��/i��8�{��j��"�̈s^PvF�!%}
�ui�&�.)�'U��U����(J#|��X��.�R s%c��>J���w��7��~��e���u�\�B��v�F�@P����R�Y^'_'�������9=�<��D��w��W�ftI:���ɬ_X��H��@4��&��Բ�mu����D'�ɪ�J��ӊh~*��o�x�/ҏ�kjD�R.<B�st��*J��@�7���5��I<DM~}�:�R;���o���+��x�N&枍�"�&�Y%=�N�bǭ����m����6������o�#y�T�5_��i�����aN`UH�EwnI�Tn��uø@�$eQ+{��v�8_�5�U��
$;�*�14��u�B�l������خ�z��q�{n�ACo޹���N�C]f�z]r/p�c��U~��h��+(	���Z�j������z��_�J��mkۋ�b�@v���{طYK�f��%�p�����5:�X�%��=��H>�Y�	���Ti4}v,�9R�-�ro6a�K��߇�&�+�x�}���Tx]4����Li�Ѷ4��L�a�* ��Ք�0n�k��׎n4�iK���O~b��{������%���j�.e�g�$�_��~��� ��&t�2_�ko�k��\(����)91����
z�_�����m�=#ɶ�S�M��&�|u:^�W��+Œ��o9�^$���˙D���)VM��قn�����j����tc�R{��'&�FH�.[������J���:���-����݋3�E;_C���:9� �LK�ZT���Uݝ<����Нae�"@;*�s���;Ͳ�cho�r �����P��r�ME�:�H���B�/�������
`#^b��J��!��m@�Z	(�6����1��Q�� [��=k���T|��{jͽ��у�8�y�#Y�uٷ/RC�U6���_��#S�������l�l�]�;^�_�-E�^�����}T���A<�X�l��V��@꬚ڨU�]�1~;�V�إQ%��_c�Qә�+(-}�
<V�~��!�/'V)ɍB�w��4A�njw1�G�&�����m䤯��@p���m *e�i�DI�e}�,:����	?�gz�O]��V5m!�cV��XjL�W_9�΅�Yc�y� �z0�,C��G�`�S�z��QNm_�Wj�4B�s�R���+b�_�WB5Lr���Ή�Ib��X�z��dYsȴ@��Lo����j5z��K~��%#r�!vê�-�� 3+W'����Yy���RD�=�;ȃ��3�}���G��O���8V�38%�F%V��4o#�s�a[�%�pDԼs��=Y򏑛��������|׊p�F�(g;B�Yf� ag:R�s{��ɽ�g`k��ަ.�:�����ŭk(]�̓H6g��vC��,�{ovH�J�뀠����ͧ���әsC�z�j�7���(�-2��O]l1i�W����ψ09ڑr4G���eP&��ê�����l��7�^ٚcg&p��5މ�}��U�qqGJU꿺U++�pb,DH���A�|��-8x\���X�ZJ����v:G~���Be����Fa�E�9�ҿ����>g�:��]�躽��Vnl�ksC�F_,d�l��މ�@$�sB8mj@piB���{����[�E�I���g�H�5����y�*^v��R�gߠؙ]%�}8�Y�p\�pr�u�&�J{Goyc�y���/߂M	|g������@5�B~��:>_��~��Dnp�L(���?����p39��?��ɂQvL�4�I��wMX/�>�0�8����O�Bt�T�tRCdG�����s;��e�B?��Ҋ�s��F�~{t�����gb�D邁�$�ƛ3%y��`�3񦬔E��*$󀠨
@M;*Kj*�}��e<��ge�[�E;�:���vй?���>8_��)@L�Iv�j�z������U��������rP����!Eўh�����k��;~I�5=��S��m�iG�æ-�7�7���ǻ%�k0�Y�W��bP���8�͞
�|B�i(Z	����]�-nA���V�����4�3"��7W)�DeM�U׻hV��eG��w�$bᯁrɭ���x�s1������4A'�c���`� Il��\-U,��å.#e��s�i� �YV�Y��BP����r;2���7�������՗�	APYHA��Q���f����޵g���P-[Q?� ��y��S�(�N6N�侇t��F9%j�Y��Ppn�B�qd<ݶ[�9@c�8mcL���Z�O1�/�ӄ���KC��I `�Wn�*����s�ǅ��h����|��9SE�Sc#���u��T�)\�1~�û��HA��&��.�V��$��a���ľx�2���bS7�~�z$⹺f�D|wh�#ƕ�h̏_�B ?ˀ΅�ڽ�x�d�5�C��S��U��O3}���S�\;f�@ٓq��;B^�¨�{
��R���鈨�(�D�)Z��5An��p�Sl'_�L^���c����L�7_p�}R��Y��j�Ȯic����؈/�\.�k�Np�#c�
1BP�Ǐq���L��3�F~F�M&��X��lQ�ܹҲ�]}Ree4�𰰗4�{�b-ׁl(g�[3»�WC�G�[�������j�(��oY����OE�՞e��.�?L����Ϛd�O�S��=���P��!�ϳ�KS��С_:�e��z��D�d�q�=�!#��
NNZ��HA�s����j|��~���cҷ��,����U�vǶTV���LC�W�Y1��z���@>��u6I#O)�Heb9�5>��P�@z)�K����&M>�X.��f>�5f�KgW%����!�x�O`�Jt��b���5��.AlL������� ӈ��4�;���YB���1��#S������0�d{	����126η�R^�U���b3TI�5"��D"��� ʝ�L�GD���e�B�_`�o���13��U��~c��@�-�)1u>:s�\�X/�y��@�>�胎W00��$�VU�Bm��}�Y�t�t�<�9G4�p�e��ьֻ����ւ-G*�U�$��jm"hx�I������lO����$ֶ����d2����G��g�r1[)�3%�~��N����HPX�/��t3����,O�H��v��wB&�5ۢ�E��w�`�w%%B�SA�@N4����@���~kn�C���g�c�
>���D8��%�WFz�2@�yN�
l�  �9\��iG�Ϥ�S�H��=L�Tlzp 4������_F[ְ㜐|�n�Թ7^���s�{���c �뢧�V7���	�̡/�R�ߟg���Y�;�o�ĉ?+�p���9I;��WE������ϖ�|P�;�!̛7#�sꁺت�0�3P���nb=�aIuiϫ�7fR;	�e�0p����/ �d�����*��O����͑U*t�J�k_+�vV�D�����3��K�5ƏS���Z*��!R��k<o%p�J�E���g��~����c��t�ç�5�$j��@�����"���� 젖R<�'h�B1����|��K����������Ev��.4D�O2+ҫ�Z�]7�$"Q@IP�)�4����	Ih��]�m�)xB%*s�G��.�=~d�����ޝ��֞O�W9}]�3'"����ꦾ����d\�O�`ċ�*�J���V��H�1�g��]�^
\�6�تy
�2t8���`/F/U��p�����sS��m�s��I�n�ϭ�H���`x�4'�=Ҋn�e�>1���A/Z���Y�#_!�9k"I}/M��|е��N>uA˩Ai����L઼�K?�0E�5):ײ�^#E��5�f�k�9����l��wS��s �