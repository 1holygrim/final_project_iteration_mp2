XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����_kۯ���rҹm�u��2�1
��c8�?��� ����(I+L��IǛ�j�f�Gf�=K�\�fqF��(�%EY�-��kK��3��&GW�.^^Ж±2X��9���{���Rf ��C�f�% ��T�o\:k�삥aӾ���~b�|��=��}�N���&�s�:�|0� ԃ-��kذ��9�ş��v�{�	*+���ѹ<2���{�$,��ȃ�%X�.]��^��V�A�]"}G�����m�{���'"�$�W\�<Q�1�\$j�Y�+/'|{[�^�3��,u����߂�f�4l{2i1�X'�
Џ��\.��Tbk��Ѭ���B�*��;5.��X���I�JyѼr[�5��!!0�v+������|c{ұC��_�QL
�	�b��G;���X�����	g��^Ƭ�N\�?�����\��0�S)LY��,���!�5�a�z�1�]�Q��ɴ���}W`����}����q��sw�S�誮����Se,xE=3o�ZV�����I�C'�
�q�]����'*t����>F��`Kᤰp�7$�~���۷~�ak���$��u�1��p����x|�_@q��>,� ���RSJ�B4�>���L!렖^�r#>��pe��E�W�j�n���$c��PڤRon/@��Z�+�Vo �ﭤ�m��C��������L-�	L�bĸ�7��U aw��B����NS�UU�k������{1� XlxVHYEB    5fea    1830@:w�:�כwL��g����ѹ��޻C�⮝��ҽ�r(�$ґ|����Nu3k���ң6a�CK�9�d��d������� ��n�&��p�~��֗��n��yBG[��I�Zֈ��"O-`.;^����D�����+�(�w;���U�l�If�*~ϴ��-����9UaL�8""�t�g@�@���s�s��o�'��;�v9}l�[��5I�h�gq��	;�R/y* ?cW�g����I���`PĞ��|k;��U�!�5�K�:�E}d�n��Ý�FL�����˰j�-�z'`b��c�+�_�"��N��.�˕�l��t6t��Q@$��������9��ᩇ�8Ħ{,�q�����#�٭ς���)��#%�3Ӱ6�]K��iF(hB��ΊP�_P�l-��u�0ĝ�8O=���yo�l��~G�z�j�̅�m�_�73�z�/���CP.�<BoJ�������!�ܱ6<�����F��@���A�Щ�x\�4i���ݾy�Q݅�^~N��6���O�R?��`㫬x���!���K�W�u}��/��ac���?�$�S�7F{Ɗv
�v�	�C��y.T����n��R�Ժ���s0~�.�,m��wpV$�9����,a���6��yPm�^N��ׇ[>n}�H#���;�4}E?e}E(�a|��R���d7/L!N~z�\��2S9�Z�Z|4ښ�ѠFxfm�@��!�P)���vvt�[Ь~�u��I3�'6��*�[u��:��Q>;Ur\�V+6�b�?��u
��޻��}��fvC%z(,5b#���U��lf�������v��	1����q`����8�w\G	�ے��(�Ӱ��j�Q��
96Yt2���l#ދrf��^�v�z1��c��Çy�/�N�D��a�p����Yvk�����f��x����O������#���Ύ��p��x��My�~�Vdj�kZ�!�l�#5|+��0л��N���uNUPn�k�7����5�M�=�m��u/����;&ЊE�rDSN�
��El��KG�WJێ���Πt��!^��5�CO{��;.|�\�I�P�4���נ�)d��"�W^�r9��V�����i������)���ѧ2��g�b`>�Em�)��9��=��Q�yG�S�>;\��;RJCl�]����6;i��ѫ��<���ȒI�5�*�堖��a�6��0�R�b\��2��E>���K���WxX7�-3��r;r��1��5F�5�7��4���S�ɓ无�
c{s�b3~�FĸG.��H} )��Z��~Y��@73�ʨ��"�Xw���O�y�K���W��x
Ӣ�kw譁��_��x�OQi(��6�������Q���Lƹ_~ĕ��2��]!�������4��ϯ�,�V�@#F���7�fU�3���:�
�z�&�N\��=T�uȸ�M�-=��h:xZ�{��m�g���Bq��-��)�r���):�θw?G��E�$И�Ȧ@x�a� �w�a�Z�6���2��<L��mg�@Y�Ί�ʕ�E�1��!��/X�3�	B���4�1�X�r���:����]v����_A�j{�+�Y���V�Z\��:QW������D����I�J���嗱��ߒ��.t�N:I�ª���+��
���C���w�L���c}��<��, <�:g��1݇�t����ftw���������vHoq]�TE��흐u��9>��Tn�9�����:�aC,Zw�ށ��nug���׫���t��F�C0(VN�jRL�r�aN������"Ԟ>]Wy�BlG�Y�l���F�>����;�ȵ�����1����ㇻ��~Qz2�GL�K0��-]�}������Td�[21�ðw�2�($d�p�fE���)!��{��Ɍ-��&����q!BJJ��5�C��=�ea�k��=JJ>�nQ�O�Eİ3	P��g���a	3�������,��h��+�E�mc�]M�x,�u�RH�T��	R�*�����=ej{�2t7?>M w�)�S���\ܶA�RY,��t�%�5�o�o����!xmx���ĕ0�1�<��8l��O�{��g���;�&�c��$04��4|�Ά�[�-��J� �"@C�˓��d�ĝiA��ՋG�}���fM�y�Q���|�y�K���ܘOY6�l����������"hR^�(]��_ |�tz�_��=ռ6��S��g���Zdg��iG+����o�i��<���X�罸� �7�l�,L�lǓ��+�Q2�{�]�}��-&�'�n�:��&�2|Y�п�v߳u����au>j��� M�tץO�l�st�� ��>6[o�F)P��z]�es�oq���~����x���'��_�,t���쪓k�S�������ǭ��;��={QZ�"�{<���g��o_ ]׻h���6߿���u��yr�����J�`��\�~�s� �j�����r���,i6���+J�nCD�����.��셕�1���y�M�w�=slz�g�
����G��-�������޴:L�4	Yi8�i/k�hF��Y��P��>SS��?$�J�B=Jc��L0�Qh�sA�e�A��;LªAh�,��Iڴl~��R�o5�"��k�E���pű~~-�Gn����T�Ne��~�R�Ql���;@�#!�gi�B�U�w��K���N��m ,�| �@�qQ�Z�<���!�cc{���ˑI~C�K�-K$��=P�}�(ŴT*e��3�3��7�@�9�߰;�z?l�+�E&������<����H���yf*��;���w����!� B�w�\�3�8��/��*Z��
%&f�S.���y3��Q��Q�����&��D�f�&!�_��e�o��_��+@�}��<����:9`�ml�B]�CO';,�&0���D 4ǃ��O=�/��5��];��2{y�#�X��e0�'j��7���]��g���v��yu��*a��,ؙ��	W�T�`<�l.ګ� ��c��2��<�d�S�T�jN�z�	�pϗ�����1 b7�S�UnL5*_��z�6h^�0�0Z�S6 \����ؠ�[S�z��OM�����ff���g5�2I�,X*0S�a�l�A�C�6u\��O�l>3^"�F�v�3��*���׶�a.Z(,�'�
����7�}�.�[��x��sm./T�9�[N���3�>/�����Dv��� ��)Y�!��M1����j�p�r����Κ'��:�(��Ky;-��v�;�m.�������#�QT+uֶ8"�11t��(-�ț�4Ai�?헺��>���Bde)֚=��a�[��)��s���*�����=SV;�϶�v��p��"`�� L������|;�2��m�w
w;�=C�ժ�*?��_d�� Ol[�LC-Xd;b�N��X-Z��}��X�}�Ǻ�#7��A�����#��x#/�I�O0�l��Ah���vڱ���9&dM�e@$��/����Y&�M�� L%�z&�8 qaJ�A��|�����c�۟�/܏��2���Wv��Ʃ���1"aP��Xs�O�H{��o�4ݑ*���9���u�WÚ�ĝ��x��U�O���ߌK>z���6����d��I�*��Dv�V���[��A�CYM�ď[W6�D���)o�T��_�Ï�{�����%3��r*�)��c,jFOX�xw5=_}f:b����,ұwlY���$���-x[PI�+���׺�t���\��A;������ܠaZ�X��㧃��8��tA����_�AE�s�Xw�Y����=�Z,���9s�Lz�&�I�}Lb�%O@��&#4�I��F�A�r���/�!���,k?�k��cUU�_t<a^�X��4[�Ɨ�;h��*��7��r�<˓� v����v=��,S���V/�h�v*�"z��1x�);!��3��ܞ��9��M����Jކ��� 4e���ʿ��Z���g��ad��B`L���1u�HFנmu}|h��+��_}U����^:<gz)lnGwZ�}]�-ã����E{�N)r�\���R(h��}�c��Е�VԚ�%d!B���M�g>_G.�A�`���$J��ٯ�� ��5��+5�iȎ�>�]��P���"��\*��Τbn�EԼd^�#���;h�
MQE��&��6�eA��Y6w>��{��k�O���?2+T��+�`;*9M%�p���Q�F�� ����Cn�%�T���Cy���w7eb%�{�[�b5�C�u�qF�z�B%o)�z_��g{���uC`�]���j	ȗX���[P<�f&�u �9�R�1婩'*%�U�K�]s�͖�Ŵ�?VTz�P�9m��z+�OSj��;\_U���d�9�s��,Q)�g&�*/��/�04O'��M�}W�;��ȕ��+P�B��D!|�4�1m������C�#G�H���HTY�,�ҧ�>*P�4�@Nr�[@��9x'q�.޳�t���c��=7	�Ake�\�G��0]n�1=�G �؟��P��{��E��-��싪��҈u?�'~��*��L��Cj�������E޴�&/ë�M�k=(Me ��b���S�Ҫ�)J\��d�ț�he�ˑ��1��X�9}�5.�t
��E1b�ć��u�C�4���D���*�p�6|�Pu�\�2�A�V��>�O`ZctI��w^$M�K���,�b���h�ڡ�Py��Pc8�/�5�xԒRL]�@��Gk���_HH3Ru Rn��`\bI�AүC��R��%���o=[I�{-aq%�RR�VP>����4�ܳ?�T�/�H%@]k��FJ-a���]oM�H]�Y޸N_|��_?{鎴�K�.��|�����!��,�#Z�>I ��\'-L_l*�1M�����"(t��J�g����eD�шd?ڀ��1	�ޘ�G���y�w��q�c�O�S�R}������&t��Ȑ�
\�,AK{�6�͐�;�� ][�M؏<�mI0S��`-����GG
p�K\�:��da�'�WSJ���[m��ԩ0 �
`	ĕU�D8�~dN\3u��|�t����T�Y��C_�{{��:�3��i��l���<����O)�ڊ�A#��ōϻ��_�;�e� t�ʉ�Hp$���R�C��77q�6㖨�����`��}|)o9_5�@R�P�ETz�,kÝ�_Mڌ�7rj��Aۗ.���j;4�\�m��u��k���|�r�]
�+ԅ�np��[:��>�X�ǳ*,M�tft�)Z2Ҥhy����W8��B'm�$�P+,1:br�$��7M|b�'�Љ͈��C��z��Z2�me4��ǐ,���1�®�>*A�qL�z�K(T��U�������b����B<�Ԥ�!=��6R��� ��@���C�_�
��G,�C����[��Zlj�vT�=��7�׋;������R���a�I����m� h�p��,r1p�(�"Q����c��� xf�];�v���A>�y��0��Jf�/�\K�)<Q 0Ⴍ�}~�tK؆*���|�y;#/o������\�!+@m�>�B����8
�L�a~�X�w,*@ƹ��3X� x?i}��'����QU�kN�4�έ����L�׃:�Ǒ��k9闄�����l!tsfxv�n�L@�9O�Jm�j���͚���ۀU���|��Z
s|e�6D�V���Z�`5�����NA[<��-�L��J�Դ&�ɸ^L�iB�=^���0�k������8=�@�a������ŇN��X�9�*��	�Ah��?�sm��ttq}������2���p�o��{��L6`���-N��{�W�L�[]��~�f����?�g^��p�Ɯ_V?�b�N�iTe�A�ټrpw��RW|]pX�%Z�����Pp0��[�����+΍���K�[���PT�S�/m�݁�}戮�� �I.c��Gj�.X#U1[��|c���t�8^�>�`*�HhxU4`a�=ٜF