XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%Ж��*�!��)�� �N�< ���n3���\,�9mk�3<�v������v���)4�숙�1v�b�fDC��<�I^�GG�q�VTЩ�9��4R�g��n	^�y���n(<8�ui�[�j`���R��b(T���g�Ӯ�̷��m9w���J��!�9��d�4�`
�KR�?!z��0n���ګ�'�W$#��FgܴZq�_�b�Ό���&C^t�S�+'́{��\Η�q�'t�{L)���>Ŋ��<��.���F��7V\hK�k������"و���EV������I�g�5���6��4�C�\3ﶵf������z�۶Tx�gί�>�����T�VGu����a�,��B�o0ͦB|c���Y��jL�gxA~���[��6���P�L��R}���˱�hVIF&�L���\��s��R�o�r�*�*S>kY���\{:j��彬X��'��P;n'�&��vB �2�jq�?�F����D�]���=un{ܓh���%�_��{Li�����%xA��mq�^��ŀv����j�"ԃ5�B�-u����-(%�O�.�籘�Ž���ew����h�ra>}^�8+�����`�з	�;�Vu��K>A
h_@ю�����{�����K�Cl�-��A�2 �UbC��)�+?����_'A��4lr����pF�S	q�Kw�&4O�)��bYS����$�e5
��z<�T� Q�k]�w�5UX^@�⏥���XlxVHYEB    67cc    1570����������5Y	�����kdy���&�B��P�e�Y�x#��#��;5kMa�B��tͨ��-�cEb���<j���uj$�8d|\a��N��S�V��x�wi����&�_3%��-��F>�Lc�b	�Q��(�K�_�<�]vI�8��!	'+l�<��Ƨ&MK��z(V5G/�#ٽ\7JX�����.9/��U0�Q��#Du�m�����7M]:�j,NL�Q�T(��g�΍�_�hx�_(|%/Kp2�+��z�ЩZth1m!��V���_,;���?\�'z��x���#�/�ٵ�·�Vhsa{�>��q	��{� �:���f��PIY�+M�qgI��h'������PH\79��3Z�������67|k�nP����uj� �� RI桓\�1+�U?�����1&N8��P�i�qK#H���E"�
���wH��ao��b����"�דs��o⠜�}����MC��  �}��������g �S��αb��z��Q�䫞`���TDL���wu�e|TOa_�G/Q��.�r�L(���؉���<p����ؔ��Eq��g"M �l��d��k�̔�C� {τA��M`3S)�1��S*�y�^+E{f�Fꟕ�q�+'Y��EX�T��Ƚɲ������j����e��̓3O�!�lԴ���Ĳ)�a������q��?��D�q�p�:,�N@�i#�9'l�����;��(�5�B�uFY0�`Ӊ�ic��+@�C����X4f9�~��QٛV|���O�a��d��{�+�a��m�Y~����X����،{�<��qD�r:��������@�ނ}q�j�sG��U�9���\G�P\�pصZU���j�z���a���u�� !`Q�.�HWV�0�.��zX�X�.$��,�r��ՐD6S Tdيc�|nv:|�|ǩI45��a�Q^XVM���S���҂�1�rR����mn�1�=���3É�������6���d=�`�8rVgۺ�bnST��(�
������W�v LlU�u��s4�{gu�
�\��z����O�ǃMFԋ��3��9��&,���1ZO:��	K�!_ױl4[��䦑���c�rM����os�8�5�=j��gFI����$Y�w�
y('�/[P�}�&�s�L��n�>��gi�]�����`�p>�a�<��K��P�g9Z�kט+*%[x����e	a�F�{���.��z^���&m��@�_�2�]�e���h�e�,;�(��ٱ�.�_%i�M�����l���=�~�c�lo���"o��FMhXg5��ԁ��@X���S{�\}��TW�D@��8���-�	%��KТ�=x���P��X�1'rW��hp�M�@�1*��w�����;��x'�Ń-gg�qNJ�kd�s�T��l�!����k�������z1S��hH)^'�� ����CN��u��~+vԁZ���ɹt������ܠ�l���V2����u���C��4K�:�vZ���W���G�]����4@�q}�qF�<�Ɨ�;�W�d�!Ρɛ��
�p�y�/��_PB� =��9��I�ެ��K�l߉)uX� F��?n���M���#�V|r��w�⥛�g��o�������v�n[��ӟD�\����;�{7Co�^���sT戰�G��^������^4_�`)ɲ������TK���)�}����̞��q��=��Ɏ��_��0"Z�#Ꚗ�W=�GOM�$_�DW3* ���C��Q��(Z�~y�ȃH��� <1�/��&�.B���r~\����/Q�(2��ia��`K֎X��0������e��mL�h��/.s��n�F�<N��\_{;=~�XC��v�3d��F	 ��v-��h�:q9�١Y�����k�8��gu��^�
��
G3��	�e��I%H���b�
����yǈ���_�.Q��E+n	s#��� $mg�3�! �f��fe���J=l��&����C�$F�%�� |�uj������xr���*V����j�g+um\�-�U��F�7�!�
�D�d
+XM/��H)���Y��&�������E+e�d��O�nK��4�B���~.���}}��wMJ� pD�/�į�]tӫ�mb�e��wW�Zצ��rO.��u��I�����l��O.�?�
��̃W���@ˢ}�[��
G[�����}$���k�"�5��lKܨ'��q�"�u���$"�wf�n��"�dmѝ��P��� �9�R�S����OwC��y��,�ٰ�F���#iD*f��.�Tl|(��:�d�)���,�χ;�88e�.����9{E�Si��SބF0�
��ှ��3�0d�,.Q��=�сY����k�	��A{Nm���4R�����Nľ<��3�=�4͇E�� !������tP�7��������l	ΡI"8;q��Dt(E�>h49n
(���/5�.����r��s=��~n>r1O���xR|��=�ZO�}���I���
S�B�E�nI[5,��K���V���a���d֫�p�T�q�4�qS`�?��Hs�i���.���c?ڞsں?8R��(�n��۽9�X���e v�(ے�{IYJ;�'6��RN~�r�,+��zĮ,��6�8�Dh�5	=3���3i�ȿ7���e`[x��#��47uO��H���B��"e�f?�3�`(;ll�_�,!�o@�#�:���g���m��9Ѹ#
��u�ܤmw��;M�oc�,�,|'�T7_��N���դ|�=�g��x�K	�n��Ph��s4�	s����
`̀�HTא���1lW*ǽ�I�����{��JZ麛I�jw23���oĮ�R4๕+5����o�0T��ڎ�A�g��ϳ῜�zEF*��Ll��WÑwr��/EV?�
a/�,�mRԅJ;� 0�-JD�}[���ٗ��ƹ��wL�˕z�����8���j_�y7Fd���פJ�]���Au�,�|�*V0}H������ʆ��;)X��E�4�z���<�#��O���˜Ү8�a��(e���I�+�D\Bv�x�&8t�������$��U0�_�E�Q�g��ѽШ��ڷ���)`��;��Ϫ��I�_V����9�@��?ק̿9���M�I�Rd6�&�Bkn�F�[Χ1F7ID?A��M�����#�+o$�ĵ�g�m���}�����,uD�^�Ҥ�<��Q�Ch�V]<'x�i�F\��  �j'o �X�~���$J��� 3�e텷�A'(:�n1�����k5`�Н�{�u
�����YY@F'bA�b�̙�?˭C��t�h�8b��k�@%0*�Ն��"h؛"%sM��H����ܝ�������)T]5۹j�\z[���k�/�M�[.�b��(�u�k<̜��j�pA�? Wwg�v� s���oliW�����`�!ڷ�����AݟB����"x7��b:~�eG�lc���(�>S2ڝ��L)"�f�Ԙ`	��}$�|4;W���6�չ�/��)qnHy�Z�f:���Kr�%l���*����V�{l�dV�Ɂ{���&3H��gJ^�L��G`�����$TT4�d��zY�� п2ѽ���k.5�q�gp�u�,�y�p���R ���(��b+�&W�L�1����6���<�
6ġ��5ڑ�Ū�~u��W7l��(�``J�vB�:3����U(�?���*����J��y���C�M�'��/��$�+_prb0p�K>�� xY$Y�OW4K�1�ep��>���r�*ٺ���p��:�A�5Y����Y�&��L6��c����]����8����"%��T�C�[�U�"Sg ����)i�=ٷ�\G�NTސ݌���B��$;�ʇ�d����S�y�K1�ĳwO{�����	�4��'2�˪	���&<��_�I��O����?��^��d��K��P$���|�}��*��f+�%��
ذ�9�~�z�S��?XI���0��hʔZ^�3��{j��D��(�
?(�r�o��������v�ߐ:�ǧ�[��h��p�������	E�h��Blcӆ�VW�������Z.��,�g�\���]ܙ��/�_[*8��aI9>^��hQ�oR(�<A����, 3!a��ǃ�jL��wj�'=_�,C"u�?{6I��c�\���.�`��L�IP��!�t{6&5A�G�'fL�E(\�=a��*�����0������HʾH�F6�RW��.t��u���Z��~m��_���{�Y�n��T��2�-��B4�������ӣ��]�_[~�Efk�#_R�P;�1?�,���t��(z�͸l�jD���ɍ��-�-Q��:���`&�x�W|��4��yݙ{z�+�]���DY��H>�<@�g��i'�K�ii�&������Ne9/��Ǟ�k���B�����*-�/>�j�~�6+�P��A�^�����ކB׏�VatX��wՄFޗ�%�����e�����E2�y��|̂e�8���oJo��?r�����LM�(�O2�����6�	r��^��C���C*Њ~�8f)�ff�$?��
)J�`\T���OC�Ru��}z����x;��cJ��ۻ?+�ZDyK��c��M����nl|4�͔�*�|��Zx!x��Y~Ӕi&��T���y�X��L0��ݢ9���$e��Q��US�����ފL����ޢX��i�*�K��&�m}�}��km�^�C�5L�ev�d��NT�?���L?d'ڪI����g)���&s�o	/�+Ds^U;��V����v�ιm��V#GI��l��9�X�U�1I4y��jv"�S�ǜ[y��i�V �W'�	Qm�=$J�í�����	���(�ģ����������P�3$x����u0�,>��?,�ūX��!�$��ujXo�6y۹6��xb�{ƥr�� ��1�&����*S�F�}Ǖ�i�.'_+�hN(-C8<��`��/v�,���w4���W.��+=z���C�� �+WɶT�c���#tZ<"ȝQ���[r�I�X|�_�Ѷ�?㤞���b�{�E��>�sxd�B	�&�8���o�D�P��ǔ��0b�A�|�7x��"�����0 �^Q�#����U����Ux�?t�j��Ð���,f�7�Rs7���S��+�Hs�A��/Z�{|�3�	F)��� E��xl2[bj͞?�����Q:i����_^O��,>&Wp�!=�k�*�
P>���b���<!�U"yEݝ�i��H��9�bνU7B��6�
7�U��:�OL	�a���2��?���B U�`��Ԧ��_V���b�R��'�k8r{;F�1H