XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��??;�dG������z^��Y��4�����jRz2)�c�r:)eB��:����e���z@��p�jR��GE�����,s�_a���J/���C� S$��k@4nx?M�
���f�zޱXTc����4O�s�9��x8'=A�����i؄ ����+�D��
v\��]�;U/��֛��[˯��N��Vs�~��#�ttډW�?���=LF��$��9�h?����m�2�����݃��&��
��N�C~��~z0�0��t�:���9�y��ἃD����� 1G�9|��V�N�Bg�Q����R �?xqҫI���'c���8�E�O�Ʃ{�NY�1e �i�ؒ�Na�����+(J}>csf�S�>�`��$��"�B��.�-�	|��{)��sP g)L�k��w/7F	��-b�e��H�*��Z�f#( ��_fw��U F���D���|�&���'S]Xjz8��e$��C�4�&�y��D��	�F�DvJ� ���a��2��9|{�_c[�<`b�jEk�Ӵ��!SF�$HP��^$�s�c�����_m�sbC��3('�\�c��h���S���"�ƺA� Г��~�Ugd�jF1����|����%���3���Zv�{�erbdR�����8 a���a=� ��������uH6ok�}Ci�ˏaW퍦�/֐4]O��3�m���f�$c���پ�9� ��N���}ױ��s%�àҰɰ��m)f� (v���8�������XlxVHYEB    a0ac    1e80�h��a�R�m��E{j��>���[b��*�����#Pњi5-_t�+|h�x'�adhčOۑ��+�d�������{�Gj�16�����ܳ����F:.L�ovO���M������K0w���D�#�g�'�`~�f`s�g�坢̓#�����5U��0 -f��/����3I�� Bm4�=aW�y޵�pX�g�L�7F�	E��͊K�#kQ^��~3���Mq��-�c3�rBb4j��X`�gl�F13�_����<kdϩ�TP��6��i�i���z�
�`�H�~b*����B�����yU�����bH�7�����������f�H$O^�Y�w��V|���������⺮��X����Qo�.�{%�OT��I�g,P����U#|ԯ��ݷ-�g��3�q�c�u�~��=ޟ����j�P7�%DoD殆��"`b:�����i�~VZ+�&#�� SD�>\,8�6��'� s�y6���"���-�.�H�-dGY�U�~1%�p�k�H�%�{9+#��ip⥹^��+�t�FNJ��J�T�䜀���5��U��"5yF��nk��!��C_tR���H�y�zRc�?���T٨ �=k�Տ�૜��s�b=��#7|n`Pp3K�mt������
K��8�}��P3���0��?��u���G�A�KϭRm_q�_�_\�6s��ўB�XaR=���������f&./f30f��	!">�"�?�w=�0 ZW?rO8�/2�����|�K^9a��Jr4�4:�JB�?P�o��Qi�lB�Q�8�n�ȃd�\�,ie�{K�\�S=�R�O�5z���qK��x#�2��*�NO�e�c'���Ħr���(���p�0hۨ�3t�g��	��Z�X��55n9�b���d�Ӆ$�Ò�B�H?G|#��a7��B�`�8�B�^��R��iA��%��_�u�X|�D{9��8i��L{s��º}RR�����۲O��{鄿���ެ��s�|��`�Sh�~I�˷"~�.j ^ȯ��	e���y�i�!tņ1������Y�$�������T-G�8��>G��r�����tu��x_�l.uq�֖0T��b�R��r����z��܎��e�/$MƔ[-�i�G6!e8�6J =ʕ2�6ԅ��f�-�}�Ǽ�: ����h��1��|�ߦ��b4��l���E�!/�y�<X%��=�#�ՌKW�Fե�x�{ѻ핛(�)�E)`4=?S�W�?s�~�ԋ&'N	�/��[S�_�w�ܨ�_��|2�͛Gd�tv�u!tO[�YU�h�o�倯�
��f���M8�E�:g�cj4�*Ӎ�%�z!�O�#駁���fP���x��7���r��E��%�{U)ʌju�&(�9�͖"&{��6*�>e��<�Qe��	Ǜ�0��;H++v�zcwF���B�E����QfAZ���0I�лE�:g�l��خ��HG��#�+R�6F�)���{��� �T{%`e"��V'�W䀜�U�N[��ң�6���O�1�.֬j�j�p�W�.4���}�t�Y�f�PJY��9��P5��2��?�K��Vh\�Bm��|^*>������nO�g*���(+�t���� ܤ�@v��/�Pa t�Fկ�u#�U/�c_&��|�rS?H����Q��K��q�LZ�=��$���C��q�������k��g�Ig�#	괯e�|�Ĕ�^]̕WՙG$���|ۮG �ЅӋ{P5�%��Q�%'R�Y}$v�*-/|A�M�(*9�g	 �=A(ki�t�1�x�J����O�ov�[���z�K����8�����p��^��wb$��:�M]�9�&�V횙��vDL�Ŝේ�/0������U-���U�jE�t�㥧&V7���x���,�Q]���@xY�凐of�~̃h�p����<7���#~,����u4�D�	��k��D#xCӘ��Ƃ)r��	G�v��5 �'���5q��gI�r�gƒ^�`�U�CF00�∉�	0;2z[��4z�$��у?��*@?'5EK�s��u�0�+��n����pƃNR*���+�S�H�|�wS6����i��U{"���z���I`a)�U՚oq�E����U�v�ȗ&${�Ŏ��!���J���6�P�U�$��@��ʙ�̑�A�9a.5(��|�W%��<"��=�낥
�R�d5����mA�D�uq����G��ҷ�O&!����Hi�����
�I��VY�D�Ⅹ*���=R�Z>9�ǣ��ϲt��N_���r��{�&����A@��
����8������������M��ڡ����H�V��fџ�D���#��M�bT���X����]>:��Z1D�������z\�L�v����}�hT�L��&��<�<dZ��G:E���4�rׇ�����T g�R�.��5�|�����I��GP�bf�LP�f�^l�$�)�����a����p�"�5V�j	����P�!�J�UՊ��s0�N!�������,b��Gq6p_n;�$N����"ػf��/�٦�]Y(4��,��P`�Ғ�7l�M�y9��<&J�����LLz��Xt�&|�fW��h� ��
6�^�W�sb��/Co(�e	�I~&�2�(�쳃�|�z�󡚳6�M��	~mС/wk�]&��n���	;
���E'{�R�{�}�{��C��.�^;�<&=���í-�`�'E�چ���<���c�.$X���t֢S5Q�V@�$*묹XJ|�e�\�˥��ݫ� ؑ���6���6�X����葽�����TV:�'�ɻY���z�Y�͜ �[���e��ʋ��y���vK��u�������=EQ��)�n�,���F4Xi��r~
T^�<��74+b{�wN�K�Ԑ��$��gP�(dW��1���N,��ED��F�7*��9�wעv(�3���Y��f��_o���y1.8P����C��L����@\%/��;��O{��;5cFq����8����ʜ�m�p�3>�>�����c�b���V�k���#�QT��Yۭ׽vD�^��Q�]�*환�֑"�Gd��Ԇ��9�1�t��kٳ��WX4tQ�o��4䪕�q��7�3���̯Y��H{F��,��b?ub!
+��tz��`ƕ ,�����&*�����<v����lD�I�1?������'^s�]�HD��>��k!_7�RlI�'~Ё��&��X�Y�٧.�Y�eS�1S$@)ƶv�G:)�����0zE0�[nM�D��I��@�sC�x���%~�k|��O�H���T)�^��� �|01W'��`Td[,��:����ni&/t��g%��甴`���5Ԏ�-f���,Zo�����Yx��1����}��oU�sQ���a]�@��7�)�è�Z%���`DN��;�_�[���O�PN<�x|N������:kV�o��tp�{���#�FO\7*���[��߭�')�yᨉ4'���O��;X����P	e�	�w5�WYpd��p�5�y��r�Y��CF�߳�2�3�ʆ{iL�v�$�Zu�I�@�o�';��Q7:�^�{4�|�*�Gܤ�,SL��N�^�K�qۂ���^��d�ۅ��/����ʉ��d�!	��
��1S�ӗ2^��ޑ�p����+\F+N <V�����e�_C·
���-����J�߈Z�[Ԁ�����.���P�
&�OB�w�K��|�c-������x:>fK�����	���^�s�R}�3��4��-�R�jG��ٌK�M�d�S+������i�5ۄ	j�i���ߥ̓�y�D��&�W5�#��iD�l�t��b}�8���!��vc�<��/Xk{FbH�t�eGd�Դ�:�2ǀ��{�>[gp���1�z��MAÄ[�,O��m�3P+����T^[���ģ�Eq��Gx�|�"���Ʀ.��ĭ��l|�^~|k����t�����8H$�.�����1Ѥ����c���O�~8ِ�"%�r@�e���\�s��ϡ,#S�=�4Q�� l�&+���g{�j4oɋ�?ǥ���ݹ��.��i"'!$O�C��.�}�] �A��2��.�#����ʉ'Q�3�������^.Z�6�CSĪ6>�ӂ��������t��X֪6�Z�m����o(�,�v?y���=z��ɰ�!l��(;�-��	�L��,X?,�g�/F��I/�x�96�Md�zȟ0g��>�.Y��Ֆ�UF;�<R�3oo�����[>A���P� F�o�&�o�YYe'yҡ�l=�����[�|����(*'/ݡ�!�@f~���*�Z*�F��,�L\�w�[L�� L���+n<�:�*��͏�9Y�F��h��LV�<���Ǫ���_]��m沟1\M�p����>�S[ ��P�;o�%370۲��u'=>������ʮ�X�+��❁������|�]@�m��ťE3i�M{����&���� ���T����l�oݻ�:,1q�=�-&Dz߼�l{����CD�kU �����9�k *�g^�bg1?�	���ՎO��F�}<�穵��!��њ}4�Љ��~(�ͻ.~1ˎ�x������4�����5��Fl��zH؝H�QM�r�^e(5�t�K�Fj#R]I$vD�MG�l�_��I]���6��N��a�螴�ͬ�Z��BGH�!�~��q�{�H�UH#9�o[j�N4S��Z��!���m�3��e0d�K��T���:��"��JhGM˦���2h�~PT�1�.�zw�lߏ�╌}[�O��sȚfG@Wu�%ac�b��t����4���?��� �QG@����v}�g���A�j?��w$�����d��Aj����Z��ϣ�gc&��q���Y�as��P�r�ܭe�x�HoOɯƚ��Jj*(�-+":�2��/ c�I )�2cqQ�N���If_�i���],-��+6 �gF ���0t��l},o2�йJy���c�?Ú�����uC�Ȼ!�liً�{�f��@5��9e��;֒I�����%������fq�,��1�eP����؉�*D�R�����zQu�QJ�E:_��W�6�+�3���D,[��
%�=;�"#ɑ�C/q[Z����c��������w��N������0ʃ��q@T��'h�u���~I���X���R����g���f�`��:��!0�Ҝ��_�b9��&�����XS6����r#-})܁�?_li�Q	�vp��g�D��5���\tL��WHb���99b�Z��-�r�y�k��rfI|��cǱT4/��g]QhSι�sXZ�[$-I�Tw��詾��F��j�Y�k������%� �O���v�&���7@��)E�?�(TrRqz3��Gԏ��9��f�$�3B���D����e,yL�˟�i;���x��E� h_:���H�?;�#
��d� ��e  dK���|���̙�y�e5/�0�pW}�o�cd�+.�{Y(,� ��kT��~W���a6��A;�M�K��YI@���X�v&5�W�a=�d�nW��M��d��]��as�(F&�HH��x�p��B�_�;��Sr6�2��28D��
k�p��<R���,��X���v��#��(R�ݫ��ڛg�(GU�q�b���\�O��>�7���}�ǘ�I�I��|���dX�X�эS\�g���$�F )�e��Z]�ƞ��������}�Q]e���	�$�a_�<DͰn_ I~a�QBT��'�>%��� =��x1L�]p&�n�/M��F#o�K��0��1E�u'�|�q�@�P��4�>*x-?o�[B�A�7�?�7u�U��,|p�i��'�Ɖ%��� ��G���[	[FJ+���E�T���䓈(0�&�N�!��!�gPI�K�����M�vO�֙E|�3�jO��F�iV*�_���c���yy�\�����B����W�ׂCu\��Gx	tAژ�8�H�gS� 73�K_R>	�t�H:Kbd�g���ܞ����Dc�W��1��$P�JgUX��f#�Ư���sgN٬B$�X��f ڞ�o�(�3]s��_s� ��q�l�G<l��?c	c��Bqv*wC�P�l֦�J5�%6L�b�2C�e��ϳ�w4����Sv�&��+�t^�f�6�ZG&2���Xז$�H
��m�{9�d��S��"ua)���X��&ħǍEY<�P����7fי�,wA����Q�U,A_
����3��㎤7��#N߮L6�!��S�՝���o�0��?TXU�J->����J�K0	v�Rt� �/����{��ѱ3u7��U�]�Z��Vc!��M���%&u*A��>�޷EX�!���<EW�Z�b��/aؽ��B�D�.k+��8����	����y8Z� %^M�n_���@�J��~���?���i�F٧}f���k{�mϿ�sړ�d�_.W̜�Y��g�>�<C��u҇sE=��߾��AH�5��d�&�/!�b�}�����ZQ�b&^�sT� ����a��2����p��ʻ9���u� �qGW�!���1#�'��K9�c{lX3��سX�7GM�&��V�R1F��f��7�uZ.����uQ��J��?W�<SI	�r8l_��

�b��4Э�p�Pн��t���vp��\M�ؤ��G��a���eΫP(�Q>3�����3��"��g-:��-���^�s��C>��y�&IT0a'?/J�1�3wGˏ*�%����{�@��*D�A�P��%c�S�3-��(P�n�?4���B��;���>AH��p{W�F��;8i��Mi����B�qMH�	��-7����/���A�l���Z�z������z��������=�K�I<b�X�EZ3�p��%w�]R�����h����8;��d�)���F��f>%Y�� �Η��6M �%B̝��yk���	[R���` m��.���Ljld��3��au]r�y�U���֧Õ�����L��E������U-e@I�y��j�?ogq���iC��/ �7�h�&@���������0u�(Ʀʽ�4Hl�XN�=j}R�v�m+
��%�4<�����N�`�ZP�i]0z��;}�
ِ�G�>D�<&0��π1�����\N����li'=vt�^W��yq�� ������1)���g̛ՙA;S@�{�$:1ȕ��r�����*�NK9��nɛ�x��`�$�/�6�&�ծ��6qH���w�dgЫ�s��^e��ԏO�t4]��'|��)�Q����֒�$�3�|F{�sB�@�b�C_���s}���P�ʷUaU��ub-���A�d���=�܌$P��#R8 ���-��W��nZ�{PQv�¼�%HU���_/�J?9�>{��:�,TTX&�[:�CR����qG�#q�A�F�뾛M����y��D����;A�Ӻ-K
O�JX�.��\n*��b�u ���3ߓT��f�8���]O�W�; ^�x�}N��L� �l���e����Ʀ����Q�[\�
ƻ�� ��!�,���S+����[U�K�h�N��:ٟ��1��M1�q�h�bE���R���