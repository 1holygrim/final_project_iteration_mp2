XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:�a����=4x��ґb���،�����8�d�/a/�Ve܂_6�H�gd�C��,�����Lh��˧�"��mf��j�*w��r0��bM�N���-,�%8 ��+���7Z�T�|*��B���zc��G�v��Ğ�����Q��w��Z�S��CX�<�q
J��g�݈`�P�CydJY�0�;�/��^�O�2�+����tA��<�FϝC�8��Q3�1b��P�Q����
)�EwR��V��eN.��Ҫ����Mܡ��˹�5'��t%7�^n�o�{K��׳Q��KT��������ռx�Q �Y�~�����N�0qw�"������,mɒ�l���Ě�^S����'O������u������C����:�3�?���bަe~�ғgf�sYn	���#d��~�����߽��nRZ��^�99����Q\%�8�	=�`.K��`�%��\^uh���S|h@R�^�U��[F���$D�G����R�X_�?Z=B�������f��? �F3�E((�{鬒�km�4o�./��HWG���S�Y��<���4믭�G/go;��InO��h�XAo�%����A�z}�sʍ'\ֺ�"�3�2%�J_}��pL��Ij-�ޯɰHZ ����@M����<�CÌn`ڪ5�`wk�_:��g��vʍ��m��,ܿ[L ��X	�+�k�����z��	,0�@e�u�F��Tu$"as���
�yXlxVHYEB    7ddb    1a30�d�S��E0�(��:�Pi�(_�3��$Ex�<�u�zn*2a���3�Z��-��'��g ���+J�C�0���~�=Y8~�'K_�H7�1� !�׿��M�M��=��9vf`kJ3|+�7�@��W�x����e��%��g����i�;��1���
Pė��(�����hGrP<�:Kh7���@�/�]j-�J>s�l�x���	N �-}h�K��	AY8f.�s����F��I�*�\`���l�-ܖ@��R�:���V��L�F(B`Z�@��6P�Mc����[��Nz�	P��L���q���0h���+jJ��U�wPWfw�]Y�%b���P8�ju	�=���B��Ƭ��R8��7m<���(;�U���i�EQ�����fZ�I�$�Yㄼ��{zœ ���yA
Zś�o���0D��j�C1�&m�F*�����d��{Q�zMRR���N�	�k��8�a�Z�Mf�/�Z
�V[��m@���3��׿��t���҂���c֖��R���A$�@�[�GA_��5iĿ��r����t=���gL��e�m��������攡��$�W]WZ�#�M��6d�z���������+K�ޅ��k����|�o:c�wt��N�o���L� 5N�˪t��m�^	s4�����MzPá�u��@d��n�#HJ���|=�,��/���R#�B!ߊM��q��⛊:�gNP���g�Q�m3ڲ��/�a�iad���B��`[�H��w��V�{L������r&�:(Z����2�xn�!�o�b�i���p{��J��|.��_�k��=��I����XA�{����;�j�u��O��?����q���iU�?ª�k���^�SCYX���4InOL�����mG{��NI>��!��ԺM���)&`�Rd�� :k��0#�z�C͝�R���4�X7��7:M�:�$�]�.�I�y���8�����7���(����?�-��#����i�P�k}�dU��xn�U��x^3�4������;�)��zdy#տ�ts^��\�$�5 ϝb�"_Z&���!�+yԨ�G�>2��De7�P�o�F6UpCF��#9tFl&>�-�� E��Y��k��%�$���_�W��\�6'L�����,��^�DҲ�X�Ub�\ƪ6A�K�M����v�Gڟ�����m��X�7'�M#k��x����,d0pF��h��mcp��O3z��uz�{�ѣ��l�2U�4�9�B�A}N�*�ҝ�T�´�ۢB��{@DA��2	�lӓ/�&�l���N�s�<����w���x`+I����լ��H�K*W����z�7nl��-���{E,� B����%ճ8��LVa%�c��w�]u��j�I=OtS�Fft�vE�v���'Z���.�j/"�ʴR�F䄿L��Yw���,`<$��7.,�h��X���-��9�L�6.>�3�"�s9��s�.�v�{֤/���OH��5�ؓ*_?�7~���
�w1	�"��)���L�	�}|"
����@6Lq+6y���y��ö�]�Z��h�b&�X�N��t�������8O-�!�z󅾁���A{*/Xr��	�5�,]h�<�i�ys-��5,��g�|�tu��\�!�����I)��e%gC��C��B�-#7����8�)��{Ch���w��o�D��'�Y�G��C �A��)��ƫ�C�q�lW�������yu�o/�r0Q��� xٛ����DK6��@�K���{�t���v!��aC���O��ew��c��+Y:~� ��� t$�F ���ꃂy�zB���h�����*�xv��N�}�,���N�9�Ψ��=�¶xr9�N	��>��,G�JY�\��p�R�\@?ٖ�BU`�Wb3;o��V�b�A$�!�:�bVg# �d���y�:ՓɁUPbf��qA��j�c��!����L���+x�&- ��,�_k��	~����kJ�z�N�98�\�[�l�rP:�	b�<�9��(��u7IeW��z�~܀8�Z׾�n��v�e=�EM��w�vV*�v�g���䦽��\�m�bE�xm�ۯ� ��t�(xx�4}��K��@��-2���b�N7m]D#+³Y&�|2e+���h5ˑ���d,�v�1��$�%�,O�UA��&��(��%��۶���r���A�G(#�n�&;nc̺_�@�.�Q����>v}C@�s"ɸ�����T]Ʊ�V��;L����>��3*�c��0a	���� c();U.��1k���>��I8ı0Ϯ9��?�O?웍l���F�3�*Q��m�J�@pLQ�(����!� �
S�������_�=�B��
���#E�h�ޫ��@��k�}��SJG�2܇ L%������郗�y����3�!ܦ!�ݫ�İׄ�J�C�~��\^�3yP^iRM=��D9�Y- tX�AJ�T�ʐl��Y������
�+��� *r!Ge�Z<��UJƼ���uԺͰQ�u]��3RxhM4�1!(iq�̕�X60�]^R)�ӻR�ba����>a�ca2�E� 95]�v9S:@C:"�q��ح+�b�!Տ���!�{5)��-L���&r�������_�w�f�{��8�vp�h5���W��b�0v�����2]��v��3Q�j��>�S��q�R8��k� �J���f�j�&�G�i&���0�	Y]Aړ��R�1��/8��^�G����[���*��gGV=����G�d0�J��>-��D�=j=����F2�z	�4�`���2�כ*�i8�b��J�d��-��)����9�����f�(&t[�C�S�7-D�<"��*�����Xn�.�H}U�U���7�nTt��5�+}]���:������jO�'��t��Բ���Fi#�[KZ$ �X���͚�t^���*hD;
M7��0Ò����� ��go�� �$��_Z"��?G��S�g�S��<���u���<UM��X��Ŋ��#��uЗ4懚~l� W�*�(��I�
.���4��P����gT�@�#dL��s>D�%�񙬈j�r	�;v��ԅ�T�'ƿ�k�v��䕢�l�(`��d�3..�N�3O�-���cS���OW6��m̟�6�zb��H���ʞ�#�h����Wd{H�p���ĕ��`lk������F��#)�[ _ʫ���1�
ٮ-vջ�\c�Ͼt�I��̍���<��o}�5)��3r8��ꏕ��{7�nbǳ�~��)�����R�ӡ��{���J=��Pd_N��Q�#����tS8}/b~Z�l��!@�+F�Rc������:%�BQ\K�����W��8�.p>.��,c	�jp釱��b0t0�<�8��o��LX,���1�.�-��j�E�j�Ԃ��S���b	/�s��ѹ���p0v�!*��^ �|J�П�څ�|���6������{��R�~�2c���Ͻ�Q��N �4�!ҽ����� &ɿ���F2��!~$����]�9]��?fAI�U�%����Uĳl�����+K�X��	��+��(£6/s��+-^8b��+Ҍ1�b��.��#%	<��a�V��K�`�d�f��a�wn\)Gn��6v�Wޖ�Ş�����c���)і����G9e����M�f��tfiWL�4���2�PȲ%L08[�n��_�+Z#��W�EV��/(hء�y�5�98��=��&9�WN�3i��c�W���k����X}8��V�m{��h�l�xSqOZ��Ϯ����|n���鮦�Z} �]!s��ވ�\�TA&�@��/��!'P���@��L� �0H����&q���"��"�Hw?S&�!PK96�*�14^�)��:՞f�ֵ���>;��4w_9���C���YZ�Nb��Z�s����GŮgwg4��Cp�(�"��])#�v0�r��mE_X��&w�|-����ydGfxT�몊�T���$D���7NDr�^�y�	�f�>���M�Q�ۅ_�Q���q����r֣v�'E9#��=�ᄉF]��l�	��]v=�dʶ�X��5��y�*P�S�W�9�Ѩ5s��m�S��'���3�		~drͬ���A Y�T$�d�D�P@��D���}-Q���h�7�k�՝��h��^�)'�^�G��gR�n�-��Mq�l
�!G_��~o��>��e�$63@��rOV1���;pkR,��*�WB�.�l��W�v�|#��E���#��;-�p��(]ȥ\�}�)=���Q lz�W+	M����
�7���:#j'��*%K�%�s�Vd��'KՈ���!��M��M�g��Q���N�J*ٱN۲F��\�~���t��B{CC��g��d�,����yS��������U�f���TN-Q[`O�s�-�������:Q��:�&W��"��p����Y�y-2���G�r����@`1��<D�/�Q��z_q7Q�<�_7H~ؾa�v�@Oו9.q-��N7չ��ѐ�?Cǟ�ۦ20~;�B�I�)�g�u���~]Ghݒ�)
7���q6p{H�i�c��<`]_�(�k�W^��V�J�A�sd����z�uR��y�F�J�IR��^�{ݹ⌫��C�m{f-��2�vǚ����N㹨?xC!s?��o�(�%����F��Dl�y�]�M�p���g�u����$��Ό�J�-�ec�|!-W
μ$f%g}@K����?��{9B�u3����h�a�?��)"�B#H7�U"��ѻ�q�*h�&�p��iE1�+�tJ�Z\�FE��Vvr�ԗ��p�n^����鷂�$�ٗ\�
�_��%��~IF4�s�;>��b	���k�Q)�/���0;�
��b�����[�w�M���$"����O�H9T��)��ܕr�l�a0��8R�����=#I�;���O�9J��TvP 'i+g�7RM��쿧�'#�mac�lCS=l��?4���򢨻��EOu*-�r��� ƠQ����G�j�����Cڥo;�x^��{`_�)dӽ.弡=�C[�So'b8�������r�f������J[��^%R1}��-�Z�ñRHeTw- �Qlj���/��jn�H }xR�i���_�}�,��yځ�� �
Xi��,���fd!#���VG����"��~�M��^��l��t���P!y�dO�\M����$!�n�~��;� �q)G�ɵ|,��k���{:2ϗe,��P��ݨ(�l�mp�˵��N�&����/������^G	Ξ�S�oi�)?5���a��6B7M����h�7tWM$���0r����^V���/�o����о���i/@�NU���w��<'��1C-,�ݘ3M�(;S=��++W�v� #I3_Ox��D���G�ɉ܆��������(�wĬҏRF�P�M�������������ݷ�L?������y�"%S2��N�ٯ��G?�(M��N�EZ��U� �|{�.Ju��l���z��ϓ2yS�w�eR�����y���/>��>q-[��9�� ����Z��/�E{��)����X<��FԃQ�q��b��-\�"�nļ�;Dl"Q����&�B1�sN��|��E�2�|������T���2��?,��(����ְ<��.���N'A_<O���~�iO�+=iR|-b��M������!{ �H�M���-���Ê��8����=z&��3�t�j���߰��6��aFV��ɍ�XH�*b]*>��td-to��uEq��J��q�C�=\3���R�u�]TγT�3	�i5��W�$���.J�72�HN���H�"��"l]�C�؄���}��	Y��'y�E�K"�%p�/��\�x�ɘ���B�t�(�ׅ_,��.��{L����EV8K,�����q.��?�#W�Q�pa Us������3���`���|�U
�!jN4��V�ݓ��~��CX��*t�s󦒱&�� ��m
��i�U&e� �6N��]@z�	t��}�����c�]�Ϫ�0��4�3���E9��+1���K3�T�Z��"��h����ṡ�0r�k�Q|������@>_��*Y�Ә�b�Ǖ��_.�H�m\=���P��ϛ������׈#��t3��~Døj�D�kF�4�'t6&L��t�Вj����,�za�|I��:�P64�5�t��8��.;�oPM�9���)��f��q	�&� ������~��4�<��1�~|����!!�s�^J��F�i�GO�xh��=��U���;A�;-gz3:P����ת����]rC�q�m
/=���|����lO-Bj!�Pf\�|/č�ǅ�t�>�����s���� Ó{�I�B�*����u����y��_�ԋlxR�L��>�]�,{�Oy��إ#�!d��/b����^�y�����w$?�'�8��>�NEBnSѶ�J%�$��􈟌�ip��ǹ�3ݔ|E�� �t���#�}	��u>��{<�t���&oiE"CoP�?�>;��ɛ�ه��