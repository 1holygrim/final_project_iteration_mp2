XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{l/zQ�����/ʇB=0�qɚk|��[h��CBg�%���>�)��^�`�";�fc��{h{dԍ��c2dT�͉d�zr�		+���
�}��Q6�i#	t�f\���[;A�r;-h����W��M��T�SXT��-3�1}�p<��I�d��I�P��j��B*"�8��M��a#+g�o��JD�I4%�p��jJ���Dl���5p��v��ׄ7�������k�=;T��_�IP�h$����	�o��Src8?^�f��(�K�T󳖋��y��������Ό��o��V�kV�s�\�ଗ��~r�=�*o�D� l>�]�OX�v�1��~�� a�r�*v��?��^S�d�����uj���H�H�${�!��fs��iBss�5jǥ��S5?�����y����lß�ws��D�a'G[�/�� �i�n�[u\�����&�Cqh���A����fyl*ƙr>ao^�5j��7��Q���yX�X����.uul���������MEvb���<���b��Cm��O���m��4��4��T]TOv�X�7�� �����պn��Y���G14�����}���L2�oI�#Z��7Z�@r��/ I���v�4<*���$�kk��۟��=���RZe���[U��ݦ p�y`�O�`���;_�E�?��m�q�[�SCdš�Ʈ��3�+ط��"����Q�X.;�k�9zPN!�ز�����I�~�Xt$�6�Ȣ}��>�}��XlxVHYEB    c804    1960ښ�#7I<t�p���ҟ3�׹�&��=��Q��߁b������O�m�>�����\��\�~Z$)��N$�Hˀ���ِE6��\.�A_K�#V<�>3�u0\��X��zfr��@I\�����5ɉ�o�R�0L.�^W����L	�>��� ��H�v�;h�\uiG����[��ˁ�������z0.y�)�e/�k�١Rp^��8F��!�LW�u�����C���J�]�-��ͮ���V�����#?pp�F��ez�~�������i�t0=X ��^(.��NO��_�� 3揫�M��y�?c��y�$�%B�+J��?����������#����1���(�0�I�y���5�t�P9<�L�����9.��>Oitߦ���mR���4�G���<!}�ԂB��{ƈ_�^ER���_S#�fx�m���W]nR8^�n%q9��N�����^�f�py��վ�!��p�ى�e��?f����~ =�APօУ�qH��k2��Q)�r^%�aCU��Jpy�[��&}��c���h�!5�t�@B��~|DxIc ���`A4k7C�"��T �����ڑ7�ֲ����~1][w>f���ޘ;�CW"Q���N��@�/'�w'xD��B�HC�o�=f���U�  �����"�`��G!+��X��N%��T�y��0���Ox2׻�?�40�J�6�5�2�}�!U���Z���������~�˳����R�.'cE^v�w����Eu�B�N��9���'x\��H8(�*)TM���HҪ�:�S\�����.p,2�̈́�	����t�!��G�y5�[���Ф�t��#A��>��VLD��s��(�r�;0�(����}�&�`"?@� �	���xeV��կ�v����0D;v����n���pE��h�G�>ʣ'DLꙧA�Py!w�7w�$f�7� �.����\@<׆N��!��T=�}��$��J�^p�Fm���+YX'LО_}�zwH��;7iZ�m 6�|i���_�U�4�� g(���D�x5J�Ҟ����IT(_;�y�V�o�
���on�_���Ε�{�s�;�/��������>����y&��o�۲9
��|A>�/�	�hJ>���7n���V�6 ��ȧO��m��aW � N!cમW���YC[�8���8�B��o��I�tr)��`<��7E�%ŠlB��u�Ž����^���&ҡ�����ap��v�O�ō�ƅ�$wo�)�9j�,�� ���lȰ)�$��Y�L�t�:k�>&�A�Oa�R��?��X	�؂y0����(j�]����C:\e�M6��vc|F�	9�h��eC��ԇmO�����Y�c#�5�)�V��Ue�d@X��u#��;ʒ�|c��(�Z��l%NF4�&�_�>�m�]c�bNo��npZ�ǿ��b���X�_�wG�3���[���9���P��� ��-@ �A˜�FJiB�����$$�z*z0^I�,f��|��ߎ�GU^iA*�q��}[����ȋ1��"��I���$�fVh��ۡ#��n-PUD {�[�T�{�|Q��V"#��~���Hr{�ȿ�,����dg.�|%i@��82ly�z}>Q,��8 2��	�B��ko�((3����h���<�*�5ew�i�>�8�J���V�n T���#�b�`�Hw渷Hl�4	��2�� ]��%A��F�-S�/(zX�D&�l޻]P�ܔ�E;�l��Do!x�$B[��9��<A��Ş�t�I�m��Cg]�Be�r,������xx�9Y�Ǣ�%�R/Á��O�pѯĄ���Z�-�"o�,Ȟ�I��d��mHPӛ�	w�z��rby������`R"L�8�@A>C@��$�/׾RKrՔgZk·w$6`����.5�=��ə��J]Kz[_�|)��Y�G�#XI�L�����H�1�n�%1����mĠb�(<	�j� ��Æ�,tH�4Ž~b{I"������B{x�-}�MEq��6ȋ��~�]�"�Q�]e��{�>��n�ϓ.J�c���-8iMH�z��k�/�4V�|��PRZŰ�A���XKwrp�(���mX��j� GDh	�XV��]vEU����WϥK�,4O�+��@�NY)����<�Zb �����;�@L8��@��s��S�b˓g.-)џ2��z��˨e����Ɂ����V�E@�`oMƒ��I��m�M5�	��GNAzt�t1E���	U"{I!�38�t�n7N3"'� "w]HFἉG��ʃ}f{&��P�b<{1�qQ���P,]U`��p|b2�E�A�l��6�s��]C[)�g�?���>���A��O��T�,�q����G�u��{��A��U���Bc��i�)�hv�D ĘK��}${6($��$�?:��y�cU&�9��=�.��7gɅG� x����V�hj�QL|c���{'��d�U	�ɥ6���l�G<�Q�XJN?��q*"8qyJany'�ᇽw�ܯ8��2B�g�#�"�;�b�:��n2p�Na���L	�PZx�k��1�-|ꚞ�̗�j.^�c&�=z��U��\�&{_!�QIT��JCL�ح����$�Y/p57d��qb�Ӎ�y#��R�^?آ������>���Уo�.�w�"z;��|�vn�wV�љDg�z�_��.���{Þ5>+���Aq�s�-�4�J�$o��M��J��w�jb|�/�Ñ �t'��� � \�Z��V���ޒ�����}vx����~������7�Pa_�b������,O����r��٥�0$����w�����{?�_1'���>�r�W�YȄ#S��y6�υ�G�O)��ZH�f�O���P= r�.���%�1E|�\��&�߲��:�q/��7Gx���6b�kw=� 7�Q����B��sea�m_�K��0e_��هx���b��`�l0G��<�:-M�W�X]�蒷�G���J�� �B�8wx����cERS��?h�S�Ѣ��E@g���q�<�˩�^�M��K����*M%1�M@'�?�k M�����4[�* ��$i͖V��@oѝ�������I.��.��b��TW*Q�f�d��8[K���*9��~G�z�Z���Z�p��q���Ԙ/�
w�"���|��>����d� �י�v\	�:�����>}�@��)s������\�D=Np�x�g�)���6��D��h�u��F�����ә~���l�P��lG��� �᱾X��l�B]Q�e��i�ovWFǄ}��x��� ,�ր�`ۀQȮ8�L����������Z��Á�I�E�[`P��@x����۽΄|#8����NF^�+���d.!�f�?k��6'���Zd���][
[ԃ5��^N'�	�z�l�x^���W"t�ٻc!1���7�����K`������>}(�;�e#�ꉕ�^M�.;�(��r��ݿ:��A��YQ��fS���+-��*�@/ʽ�ܗ�L�)ǩ!�7 ʜ��ʗ<j{��O\�h���߄��b�`����!���ޯY��NG����e�h�������~<�^`���U�)x��X��-����0�U ���T�?6).�U��Wj;�	Y!�R'���p���5�c}�1���qD�孞�i�����ڨ#�(�(:��ڀ顣��`=Q�,�_	@�q���z���k��@���sX�����K���G�Co�i� sfm�
+�8����J]�AԲ�u���d���8�}a4,}���*��cE�%����%����@�(*g䩮~���4=�pUG$������"�Ÿ�/rW�??b/ڇF+�%8:���h�������}]�ڽ��O�X{��?7fx(��O$�|��J/�Q�t�9���?�F�:���]���r�a_|���­bd<�/�3��hCn^�&Ⱘ)�$����<��%�����r�ŕw��O�΀\\
�~3���c�`U�s�0���cP�Xw�6�]���S��eޮ�e{E��H�+e= ��'����r��M��g���}v��v̰��nXExg k��>���.1_��:��u����������l1syN�{v%�Hu
..�R�?M,m ;P��نQm���|��j�U���Va��bSAw$�F�8oy�j:�(a.��t��¥��]���Z:����+�b>�r���SYL>E�	�K�f��w���;�SN��{2�
k�>���� (A�sTew�X����	��1K��M�����ws�e5E��n�e��q��^����zK�͂"�h��i��s��j6�7B'�����k"Q��q�� ������r�IG�&��Ȅ'eCQ��e>E�J���+�����>�":"�y�"*�-���:����l��v�bG!"�>m��>��.f&j:I�@ak}�M3��s_�E�_oނ�������.M6(%b�Pq�&�榪��["��U���R�%_9�M"��ݠoY���G�&:��P��j,�����s��*������b�n8	WŔ�)�ϸ�_q���#2~��D���9���d�3MdǮ�Y�P��;����kІE�c��h�"<�,�J�q���l2$��b���m�	��'�(��Ia��p��&��a_|���+��w1��SYךÅ�&�w��`%��w��3g�!;E���!����v&νhݶq�y~��F�}�b�e��Mh5�.�]Q����&���hm 'x�ƽ�_HR0>��-�Ș�q(&�C8�(���KYa�ꅉ'iHk$������=���G��v�i9�֣6�}Q�M��I�#N,�2��G3�41�G^���^�� �VCm�oi>V$��Flob�l(��|V]@Bd�c��/���;h��������?}F��������G4�uh;pb@ žjLeW`K"Dw�.R��1��|۷n�>q;�A�����*Su�eH�-p���%vû�2/Fn��Ʈ����~����í��(����3r �ߝ�s>�S/��k,�*�E�oj7vة���s��adz��@,aT��)h2������臷:[M��v�'���M�f@[��R,��H:Y�ʵ	c*sH�>�0a[~�vx�SL����A�k�c�3���\�a(F}}�Lj�lj/�Ȃ���6�(gL��o>�4���ݨޅ���gUu�Z&�6��Ne�Tj��<�!X�#bP�����h�å
��Ok:��w0����u<�]��|� �2f=���E*Ps�WD�:���@3��2wA�.m�d��,�u�W��|�6��Y����Yk����t�5v5�n{��=��^3�����H��!�\���|�l_V��K�?����p�2Λ����#QBو��B��:��TI����h?6�A�&IZ�P?��8x���z��B)���8Ѿ����5shZ�D��)�7�a.�_Nr1�CX��g`4s-CN���Q�Q 	˓�:�.`�!-Tc)KFFB���D0;�����C��W�P��GS����vP���Q��'i�sIǶL�S�V
 �y�J���aR�
+����������������d�(����]2%{���t�[l����w�P���5�$���'Ӏ��Kjt�7�OI{�Ds�s��du���������� ��C&Q�j:i_	��sw�<;���L���9�8P��[RS�@�>�̔ೊ���wI ]�Nι��`],��~���w9�H���cl�dq;�/����=OX|Y�
\�d�|e	��e�s��[ri`�-��9׶58�X@���M�͕��P�6GH�����!�'�P�	��z���Z=���Np/.ۊ�\�8e�z� ����)�K��&�#ҊhB-�͘��5z�(�ݭ�:$KE?BA�{��P�� ��w��^$�>#���-��O�w����u߸M�N�6}��_�T�>�hn�[� ��}�ڱ�������YQIʑ^[�h2������`S����nƞ��ƻ�6}N�'.��6_�s�������f��h��jNr!�-ٚ<�]8ȬMv^Q���}��\�ht�mv�S�0{M��~0�WÝ
$4��R�$��ߴ=.YӸ�i���F?N)���I��i��M��$�e2}7!H&�=L��Ue#�re�D<
�vg��Jw���	njD ���両w����\!����Z���q���8Tq=7�i���?�0���Fn�b��Y7�)���v��b�E3@���LA�D3� �Ly�uS_��a&�Z�l=�fh�l���K�s�Wc��(l�4�|q2kh�