XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c!n&R��,h����=��E�b0�I�'W��c��JaA�+"Ao��4�'��]/Z)�����v'[��\��a8��x�M�	"Ĵ2I�����A���l�j��<�h^�s�D�b����w5���V2��7�
��^�[�z�K��8 a�d5��5�w�	�+�x�A_X���[�Y8W�{�~�Q:�P���z!D�X�	�����vJ8��il	_l(���o�X�`����?!u�23:%���+�h�ڷvX�k�����s�f\l����e3�8�Z�(����/�]�&W\jh�ޕb��a+a$�cťϥ�*���jZ7�J� ``�Ć�%���ώ]	k�ˈ;��3Y%������Tw�j3�Y��Vz�I�r�R���Z� ���W�h��������	?�F�F�ܻ��l��83�3�zP�Y���X�M�`僮���K��V*.�*R(4�y�\�䄅HA8�Ԃ��`�_��0*�"\���_ZsI2)@�*�C����m �v�	��2�?�����A�3,�i�uG�n�i����o��V���7B�u���a7��I,P���rzQl�?{s����W|T\gx��V+����d�>�`Gu�W��gZ��$m�A�%�vO��E �d�ߓ�F��ddɬ�Lr9��;�1����;��sؾB�T���Zp`2E��=�E���fD�օ�E�#>�9^)7�R�DJre�ӆ2����*�ݤᲧ"����n��Ҝֱ�׍K�ޘk�|$�?�����b�G2HF��XlxVHYEB    729a    1770vr@c�C�z��a'OYD��ͷ���8V�m݇�v�z�ai��n����?�3������_܂��	��i�����[���c���`6�o�i��χ�u!S����w�BC�Z��@L���1��%�Xҗ�x���g��D?���?���	?�W|���;�\� MAw�Z�P�j6�cp��*\}��ş����w)��B2͏{�%b�pa��>��Tҋkz? @�	�q��Ϛ}f�8��w���i0��\!�3;��u�I��TJ%��=���^��o�zVҔN�_�;�tp��_�7���l&����sO����я0;��ޅ�ڰC@�l�|���>jz��gY�K@�U��X�/����Oώ�Nn�@�����ڦn졑!W������u@��lg��4)##���W?0d�VPy#2����l�Ҩ��hz���TT4h(�04�B��q�ˮ�e�A�1��/�2�O��M�����Q�q��/��F��u����|s���Y�[31��@�;}O��r*�����VAdT�N�=U�?	%[�E��щ>{]�k� �05�k��4C�|I��)R�3_����z)�l>)��[~>��2*���O��C��L/o(Q	9�-\��"Lnt�
�HG��Un��Ԑa6�+N,�r�cn8��EC}V1����� d+z�&��>��n�Ԭ�Vͤv��T8=�Q�7
v�����D�b��~/1��O��#��٦^�Oz���ǗbG��s���R�~�H*KƯ�o��	�{���c>yG�y�M�
tm��J�'����e؟go�B��
z��9�Z��d�yA�`������݀���)���g7��'x.��a�/�24����_�H.����x�H)���d��X�=K[
G���i9Z%-V�a4���ȂW^�`aU� E�M��X���y�;��q��"��[X����B�k��n��j��02�x�n���Je=#����4&�g��9���֚.� �h�@����h�KIt#��-KK|W2�,Z_ [\=qy�/P�+� Y�,$_+�.�j �W���R��|�RRӱ%.��������1uȎ�}���?�r�Pa���(�Z�&�"��ȥ�m`�E�U�B���?6�ՙ0�SIY�J��oi�F`kYs�w.����'�Z)&� e�ם��8��?���s��h}�W�6��`D�r��N��߹*:���3[�6�j����y�W���h/�{x+h_��γ㖾*��	\��:�=�<+�s��y&���A�˳.'D��t��<��S�����ץ�9�X:�M�W���k﵈�
+rC��C��8"�x�bq�3t؞����ѭ�SY���g���*���%gzJ���l��M/MmY,�3zݜG����2�^k8	�y�s�����s�P;���)Ԧ�T�=t��+�d��Fy�M�ڠ(L�H���W������y��^�$'ff¬�/o�}ܫ�Aљ���.(��,t���n�KߟE�D���8܍M�F~�18�J�v��)�A�^�F��+g��Zٙ܋�ã'�����Q����5D�"R��x�W-5���V�G�ć��^�`��*P�C{O��G82�ŏ=�e��iG�=�Sz"(7��ٻ�X]�%�2b�~հDrg=�E��
4�'�'���ʞ��U&mG�s\w�;푔P<����Q��ku�f˭[���"FN�U�Ʈhn���+���e��B��xoU�fT�R�����l�~0˵��ۄ��\���Ż.z׫�\���k�� �j�39��Q���EՒ7o{	0�Km��EO�6���`�t�/�YF�#���z֗��ٗ��"�UO�rϼ�V/ͬ�~��i��f��@w�n�9�Tx򘉒{J�ԟ�+������@��I ���W�H�.	�ӵ�9z�4�`�|W�逥��[�Cb(ʘ��l"�B�3d��8=#jZk����I4	7`3Zc����E���f�ZlC/֐=ݛ�k_�|���J}�-�Q 5P&"�4�66�2���[�;��/��_�khoyy@cҼp-�WI����=Q�1�iՓb?��CV��j"����P�G�X��d����ަ'@�3�a9�΄���c�{r���?%?�+}ڂQ���\� !R����9䅶u���j�cb�!�Dn�����i�U��Hh�_�q��,;Eo.Z�̻��|���8b`��s�Op-2#Nd�z�P�FVM���m�o?|����ی�DkB�O��'Ti���\^�9
�L��i��Oac�~��Bj;f:ac�g�����[KI �M$�oN_���ܽuĊz2��%�ui�䯀��<���x�ݡ�u��E���*J��s�~ڬ ��S��ku��XK"%g f���[� /]��L1�ڦ1pV����>I�K�b��\����"�1~�t���q�g�w,]�H5�����f��;΄yj����̥"�En��f��UU^?-����MW�[!X����z|�N�������br�P�Q��!�Q� J�G�1��
�svѢ�ep1�x��ntw;<Eۣ�׭�[���|n�)O��&�ɹ7�� |�Ѐ�+P�� i��kQ(Q��?��_ݚJϊ�D���AB��Ʈ1|/���<:������l��hI��W��s3�dW��Q/�.�~Ĩ%nS4n�)�G�K�z�bȁ�P�mⰇ�w�կI���U�+���N�������(�����\l|�a$Ov>�� ����J�ƨ��H7*4��ytJn��{�3��C���U�f�J��gd�7ʜ��'�|������Y\If��P{�����8K��̏���1���r�o�z��
򙁮B�3eQ��r�ѷc�P�|�<U�(�9�.+�k���ٮ��z���T#��lQ/�Ęl��f��Z_@?_d��=�>g�p<;��d�#�fȂ��<�;����csў��h���*����m0'̖{�H�6�� qx�B���V�,�d~,	3
S��K<ib�b�-�+�P�Vt�W�J�@�6�۸�u����1��I�S{�Ч�<B�T=Y�v�J08��s!3��Y)t�t�}�s�a,>��f��;X�͹��"��f{�C=Ҝ���i9Op�8�f?��ߣ�p�D�'�6`��M������29�S�ϖu~��b�IA��F���`�{c��/��h|�"-|j���zx߻�F_	"�hJj��&�r�z�n^+���E���P̎��/��R]��t�!���1���^��~ngh.�a�Q��#j���m (�N�aQAtHq���{ &��+}�"��W��nX������#���~<W�2����l��Y��N�϶u�Y2�1��A�Vl���:�]���:�rj[�����A��RU\3��j;mֆ�����t��Ki�����2������^N�m)���{#��x�rݬ�en+#�����May�N�`ƞ��ѓ�>o:�X�P����U����܊V�W�ڔ�.\��5(�f(c+c�Q�E�%�'}H-t譛��˾���پCy��![���+���=��p���"'_��ПI����}�b����<.�Qt�V=e6� ��a��H+U�U�ލy�T��n��:�P�$����v��?���pM�:2O�����ɯ�ћ�z�j��N�"ⴧ�&2o(����wv;�O������[�x��&��L�v��X�M��H� h%��;ą=⒕B�<�'�O��+�%`���*���()q�-2�ww��˓�S��큡 �)#Ǜ��F�C7�������6ƌ��j����zy1j��b�0��D�erV��0<�J�y��O���\�K\��Ċ������A�IHd�j�/73��.�K<�a���r����i��Ǔ��>�`L�ȖNC}�z��U��)5�%w�7ʛ�d�4��/���\�T�y��(���s�mDD�|�6#*Ų��'G��W�� �j��mV�u@D���Gvm�z�'��������#��'õEf��5����&x��3�]@f���B7�X��G2L��O<�Eڠ����f�c�y�k�7����,n)��>bsl�qMo"��ɚ�|9����pxD\X������{��1��pr-Ӟ��4I�	rT-B�
��I�i��X�@��ך76�~>���>�B��V�1�A���7*�ñ���s�6W�8vlBr�خ�W�����*"�A~W.��=�-��Q���t��3�=\�oxC��N�e�͈�=��n��[p��>%ri3�F3e�>���r&
r4�<��έ�&����6�eL"7ӷb�Fݕ�����P�D���ym�R���m]�9�b�Db&���3�3�L^�+u�����խw)Mzt`��!��d�S]�,ԼD�.���g��zЋ��ώĺ:�j��M��ΰ���K��CTN�@G�M��>]���KJ��U�fU%,P<z��	�5��%4`�	���B]�e��>J��*���� e	u��\���]�Ϧ�d;��b ��B����4f9n'7�w�b��*s���}婅w��d���J�rg�u?ȳD5�U�y��r˼��E��R�K�D�.�%�s���f�M�̆�q�e��s�yĞ�"��ޠ�1Y�rb�]�)�O�!@D�I�N�4��(��/��ڕ���o�N%͟.�&B�r�q��	�{qN�2��_�*�=�����������G�N��o�����P3� ��@�&�x mb}��r�_��	z]�A�DD�D D@�ţ�Ė�B���R�o�^\����H��1yd.S�A7k���w������Q�?�1�Q  �|�}�ΙJL����_����œ�y��TAh�i��cH'ŀ�c<�2��B�=�6]S�Ҭ�HuӠn^TG�� ��G/6�a�{�G��p�N&�S|Э;B���/�����"�N#(@�[��ǔt>^�V�Y�2�u�|��&$2*C�C+�d:VV��g��	��V �葩�'�I$�`R�m�N	�keӧ�`�e���z�ـ���}"x���%���*��N��ҕ����X��`���R�dX!'"=滴��RP[Z��Le�\떑�3�6�O���˨�z�Q�S]�����Z���* ]e�������/z�]�R���j��L��a��S;�=5�w>AH�>��ϭ �`!��b&-��>��-�4+�q���_�bUmV?�R<U)�-�"8�)�H|�.���Yx��>�M����#`�Dүcl�~���Eۯ}�/W� S򱆽��U��5z�ؿ�(�+�E� i3J��}]��M|��	)3ǜ���[��.��`r*5� ���vp(��\�f�'v��mʟ�/�HB�m@<'�Ŋ���ɲ��7�A1���O`dt�����|I��������1��(�����$<�ޫ��p3c�5X垙��3/}.vk'����w̯y�_��#��'e���Z��m�y"r/?D�p�ӳ�,S�6ފ��
xw���-��W2��Z0��~\a6����=Z ^��������s��e���K-Ք���]v|h�c�(�ף��&~}1��g��_���i��A �-(Qh�[y���[8�ɤ�k_`���9�Yۻۥ�(@��i�{�R@ ��@�e��-T=�9?��}�n���*�(�A>]����K�p(�����7Ϧ�Y���}�W�x��c��f����s-�/�d╯��q�%�*����L���}ը�{��af��Rv����UN~@{�"����"�ބ��{�+���%Y�$�#�	�Y)�('�Iޒ���'j�Q���^D�Ը��b�~�`���8;��r���|�+�~�;E��