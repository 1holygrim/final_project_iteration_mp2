XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1����p���:Ove��7o�����6v�OEH���t� Oe��8�*� ����'���?�,�	�(V�˘*S�v����Q���i���-�J�$5o6�ՎSf	���ؿM�6]f���D�{;��<�`U�Z������������x�;h�@|��~�w�K�B,ϫ�Y{"�?P�B��tE�� )�j�ly�����>dr�m��0�m�Yτq�qtj��`�>k'�_bΑQ��.��el��
Դ�����պ�u����Z�݄w�}����2t�+��[�f�B]4����i�kY���R�&@槎<�(���8�ӏ���P����K�0v����U�S��tr*
x�^ǿ�6��%��]
�!w`�  ��4]�gFC����<o��KEi\N#>	r~�zRBd�5���
>�!|��� ��A��$�������9�����>����6��̃��5���B�:��T�2�kd@{�����:�R��xS�	8�#G���L���A��ȡ0l��Q�E� �^�繵"��+Q҅��&�~^S�_���@L҃�G�n9{� ���l��h-���l+�E\��_��I��V�/��VW�#�S��;S ���T���^��EuF��x:�c���,q��^�a�ՠ��!�k�G$��2B{C�[}$CDP�+��M~N��\LH�&d�𜠰��>��4\\� ��W��>4$���E���a��u!־�w��6ys(L�X�(�Mk|BXlxVHYEB    3b09     f80$�.���h������M�'�	��aRr��L�Z�+0���L7����x�ʳ#�FI�f�A��jg�$��<D�K��(s���}zqLt&Y�֠O�HS��/���k1~&˹�L6�
>Vza��5���Q q�!���f������o�\\�y��
eT-�wI H�պ~�ʄ@���0�Sݿ�"(�����2���V�8��h�c����;�N�d��祛Oм�l�}�ն����V��5a9r9�iᏙ����
��{������xk�����1�l��Od&qB�C}��cݓ��*v�1�gi��G��rdq߮!���(-�R�J�!�.T����JK!m���nO/��C�­C����"C?�C�&�"��W��|��^�3�J�fu��k0��eF ��=����:{Yiξ�U�;��~)����Jip�T���ČK�X��"2�,l��6� �$׆J����,��ݮ(�u��c!@ǀb,�i�#9GXy/)�P^ZF�6��H��<�ت@127���/ҙ*�@ǎ�q�&\���E�t���tPL��[\���ms��q��5i��:|w���;�e7���k3N2���.`�8�s��ҝ�ߍ/�r�z`z��J�����3T�K�����$3W|6$��P��F}`�-OC���}O�XƷ8�����҅�*w�cK�e���W� -;�l���Ȳʛ�\
�1�ȼ(�	���l���p�MK���\�V�q|�|
 �������0����9��f.��6|֊U�*���_ǈ���~A{�-��L6�G��ed��ky:S���7N�/�&�M�;�z�b'A�	&���v��<���?��&ڱ��Ñ��b����"���\6 w�2[���/as]�4�����t��g:�~h�@���!���{�3�t��� �}@��sF�	�^w�.gK:k)�\�$d�������+ X��@��p���f�-֐mQ�x��+ы��@3�?m<�MB��zR�y��P\%���$5>[T~7�	.q�����@2k�̵��(���;�ݗ�?>��$� ����@sm�s�J���e�x���10e̞��#UX��F��zT��:C���ې{S-%��=^�7���L�%�ͷaŘ�p��<3�Jj����D�εO;��~����ќ%A�7/����s���{����]�!�6�F8 �=�2ӛI�2�q�舌~
�ϑGhi�h�Гgt>إ�?�sJ�x�R);+����?6ۙ^Ka�g���^�ͷ��D���Tr�6���.c����������O�������ob2Ut�?7 ��1�Zcn�OF�����*�������q����&@�������Y_��'j��W�|
�t�R~;r�p�و@yn|W�\�Ν��t��r>�����T���$)8����G�cC�<�f�<����Á��d1$��+C �=g�Ftq�>��*R^����IV��m}5�y���0��-i��c}#6��B��7_��E	��A_�;afa�P��>T�az�����H�x��\݊��u%�/����z0b@#��߅p��d�o����HL�h�rN]5t�C^m��Zc����Mu�l��X��qz��%�V���8�5zyM'�7��+ljnGp�?2yt���_[����3��ҳ�jK4\��d���`�(�jIl� Ƶ��d�Pܼ�)��)�(ٹ�&��Ɲя�曾pޱr[X��Iү?*sP�}d�T<�5�t�پ����zN�j< O��΢���?�zÐ��C5���B���)TB��o��c2��Iq��<ܳ�,����< �w����+k�->W ���L�$Ϛ�Z��;�c�/R�#�;��?1CE��_js�gе��2u�����"^?�>�gl2�|]�R�>4WS"�VJ,���yp�Cm�Wh%m� ���L�)O�DW7��	0�����Ɋ�y�<�%vAQ���w��Z�CUU8g�K������0ogm+S�3Yd�]��nuk�0�ѢW]s��Tf����K����DcҨ���$��Q3QT��<���\�5V(u4�x�g��;ͱ��^,��r�0�\�qE-M^��h,��tT��@mC��?�g�����k�u7g��xL���kd�aBP��ܢ~�p��W�EL�$�=����$ͮ�F��]j�]Eh��+�{�q�ǰ�q�T:�4��9�I;=a��*��_�A�V�'�y���^���LTM/��,��`o�O8��B*�4(B,�j�=������X�ؙ��
K�8	���TԿ�.e������0�W2K�6�E�j��ۣa�E���]��� �j��2^O�2�.����h��F�ȝ׿PnW��@&D�k���)���4��,������o���'Jd(T���b{��f�g���K
N��o�K;�"�T��yaHoC�[pƲ1��(.���3�E�ܒa^�յ�׬u���//�q<�!3�1�ժ��(G�
�	�{��}X��5�^�2�'���GA8K��� ���WK�0�5kE],��\�9��0+CH�tD�����d��~5Y�仼O��-j�՘+F⭚K��{/0d��5x5#�s=�#��q�/}�"h��oī����<P����Q�ڽbTxJ�	�H�4�������*	�WE,�5�Y��1u�D^F�gϿ<�Z�r��
���L�/q:>sE��H�Ks,8��t�)����&�_䦗�}�Y�|�I�N~�z��f�ؓv��xUVklnm������Á9ꒃ���i���+�5ʴ�$ax��h�}����g@�P���>��)�c�u��5�9�Q��ϦJ�r���y�zU>�+�
÷+Y��N/�~�P�-�or5����@��;�X��^�%��!���_$�%��jQw`tʙi�s�Xd�$5�c�)H��j�g��)��U���gf;<0�v�<�^��A/#�܆��-F��N�]Vp��ƭ�an�f�iɚ$�Sox��
��J,k�mt��-T$�p�!�j3U'��1Ǎf��QR�p Z'߉�tz[EKM�xV�g�r��Ə+cl($,A�����{����ma-҆�z���D���d�_ڥ%,I������Q��]�c��p9�b�B]e�Ob���ya���i��LL���ѹX�	�#=T���tbK@(���֒�룜�Gx�QCU7��ͼ2X���{�iD)L�܋╄j�#�:K�e�ɱ���1�~1l7��	O+���3�B+`�Yb�Ȱ�p�/ε�#֞.	�V�I��$ʈ�*�|-���d�������	
�*uᖵ5m�k&����ζ�jnp��ԹW bL��?�K���ׂ^��-`=Z[�K�	�C��%<,��`T���`s�$�i����=/��bbȅVS����(�?4�6Z�,�t�- u
i�F��˺�P�"�T}���;vN���񘟔�ѱ 3h�s����D�d��d΅�D_%+�Y�o�ЋBk3s.��x�Uêj� ���r/��q�h-P�r9�ri_o��S*�t.~�~��Fh��d4�<]	�߁��,�u4^AQH7�����62z�����p�n������K���N��bv6x�ܕ`�I�XG�e�$��jK҈�	&�����퓵s"��>]Ӧ���+0�{�_�]��T�:>-�G>�y�yURu��WW%� lO@zrߋK	�|��I���1L�p��A܌�������e>k$J�p�F.S��N?����w8��}g|�+�Q^gL�X���M����ѱ*�'�-��w����9�/�.��ɏ{5yM�P�7S�e-%���q*IM�J��ye`��37{�I3���k߭�e	@2dO2O5s��B���k�Q�EF>�uS؜i�|7