XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9c��&�dm��;Y<�E$�0��>��:W�Mwc�t��l�M�_�o�%���B6ʖ�����]A}��KՋI� &J���-ٜH{-*N�� ���ܳ9�48����a��d9̯�%�E�c9F��i����Do�"�.��!q'��\x-�%�">��>�pI���V�2���a������0:�e�O_X>G�+w�tP��J�%�t5��h$Z���~�a~�#��Df�k�ezN�A<�%�8%���^J� AK�9/+����j�4�x��;���q��l<q6�" ƕ�� ��U�v,҄�J�?(?��λ���H�|WH��e� Z��� ��� v΋�j�g�In<l�ˇ��������������5f+Ο�X!@��|ju�I��2U�Z�����T8�.V^ʝ�x�i&��B��������gVh���3K�����*�W�?�]��.��x($IǀX�c�8Ju�ʧtr9�}v��� ۳�K��u#e��y�ц���(��x�I���G�%�ޗ	H�X���R�ة�$0JC�Q�3���/[q)����q�83*5JI�_���ޅ��+��x<�[ή��⨑�V+�O�|��H���զ؞Ǆ��c=t~ۊ��,����OE��g�:�T��`�Ò��<���.��%��k�8j�8=�MA&"�a�eDa��J.c���{ ��wN+k1�:Ʉ(:ZR������2�?���3��qg,K�9���j�\؊'��낣�G�XlxVHYEB    2ece     b70ȫ���6�r~X^]��w�}������]��-�|M�Ӥ����C��9�C��n��TJ�տ4,�I�M=�����I�Ѫ�r��8�&N�%�9�y@ԥ
R�����{+&&��O�XTGi�ӹo%,j�i��SAq�}����l���t�@�T"�f��=%�]�n��L����.�Ɉ��g�(��W�GF�8�Q�M4���瞝أ�i&hq���ec�C�����~ۃ���,��e೔�L�w͖kH��cE�u���)�$��f���nPk}�ea�	�RwAi�ߘ�m��gy��!N�Ss��TA���x0���0��ә��Ѫ�g[�%'��'�&� ���ӻ�� �#��Y"�I>.41��#Kq@	حs �E8I�S&��ϑ�\s��*��O��ڲ��8�?=x+��c�fJ���XIu^�k/sW~5���N�ŗf+���ҵ~�:d:��D���8���GϺ�,��hI{���|e�e�K�.ٳ7�t�T���P�҆������Q�"���`^��)��q�K�0�����|׺C���)�K�t��*�>�Cl��#63��W�_���lL�Ǡ�W&��P1�	���/�9 �#�ʰx��'��>D7��BQ�M��[
����`����@�TVSAm�����qh����v��\��BD\�)����P�`��_�\/�<���l�;Yj� ���)��S�EwA�\r/����M�5�9�K�&X���\q���
�*����sՑ�L�i�&{28d+���vej��),��Ɲ_'��[v��_��8�$ ���y�v�8�p�cl����<�7+�Q�m~+��X�߃�G2Ϡ��p� ;ş�C�&h�W��|�}�����0/%N+m��\�YE5�^\��'s	�:xu	�;�F��G��-�T!���UH�
jw��OVEm��9�
�i��t������Th���0��Ŏ/�w��j�r.�V��e���gV���9+~�ה3&(\��d���R�0^���3«�	���F�o�!�����	�i-}'5��C���3��-(Z�UgWPӪ���n��5,���Q(��ָBѰ�0��eλ��������t^'�?(;Iį0.�T	��\Btn�f	>[�H����}��0K��U���ՠj�����z�{�U*ԗ����@��%�����+�ҥT��We���Du)@��?��Tn��iS�j��b�RyͲXt����M����2W�9�cF��J�1�� �8�ßaqW��I�,�G$x���V
Py�C��L����{`�cI���.�������)�`���"ThI�p�r:'��pv;��p�QZY}ս:Q�b跐�8�8�O�!96u=Sfд��?�K�"7��}̏��r9�c;ٴ`S`�͈��� ;�.���K�V�B�5����@hk%�dL�rQ~(D�^Z���׾�-��M�}+�r\�¯��THg���F.�79�ٯ[�K��Wx$�����C�����m9��:��:���+�<�p�u�k�q������u ��u����ɱR<$��k�d��*r�v�$�:y�C�,-�9+�Yٯ�rނ�26��K�����k�*�h#�|�'p-w鲳Wn��3�>��t�=�5+��0%0yع#/��qN�C�z%��5���``��"u���n�CT>
�?O2����7�u�>�}O1F�L�↼I.
��@�w�>�[\_ �bC���ȡ6��)1#��+��S���tV�;U���Cs��Ϻ:25�;�po��b�H��*�W�l@�]���Â�˩l^�	������D}L߭o�tu�K�}8*6Z%)u^�s	���+!�t<h��]��썹�O�F���X�������=5AP����e�8[��)��d��+�&�W��T:�&����d荕૒e�6���-k�5 
�T��X}�}V��Y�&D��.ph�[��wM֖�������� @ı�6@�tԘb�k�qǞ���0�\��N2?p=����b��ܲ>+�H��%@����7)\[+3 I�}�f�s���M{�ew���ڵ�
.��k`%z���kK�Uu)�0j�yRE�n|�
k����,k�}��b%G�F�<�֬D����-������Q�<��'1����tЪ'�nu��a��h�(
���!��l�f�����Y�o@�.6v��"E�D�6	EB.E��ơ{���������<6��B����.�G��/�7��#�x�,1��j�7� �Q��y��<�g�� �>a��TV(%٠m_�[�(}E���)�Em�-��m���K7��I͟�0��W����/ ���}�����B�G���w�YLբ���0m�_�����(��}W�;�`�3��� �Bup`��)�~�2_,���Wn�,�F<��^�'e�8E<�ӟdp`�e��0���A�[��0���AI�x��y���H��C������[��uE�<C�ϴ:��N��5]o����O0:ߤ�K�k�A���1�C�Sj��\�P������DH���Z�  �{�����b��N��n���h�ۥ�IHZi�Fz�lm�����}!�Պ݆���y��Bd��4��̀��c�������*�q���Zo��w�"�H�u߫�JO��.X�k4} d�1#~���̚%���HF9�u� 	���2tS�'<@�g�6�ƆR}���m�'!�Q�z#���]��!��)��|�!��$����ܾ3��<��:q;��+�������D��:��֭���j�������9~���ʙ��fC��V'F���M�	Y2i濯�x+y�Z��_i����栂�[633�"�Xü