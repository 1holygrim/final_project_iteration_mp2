XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����F��ݢ3hN\��aڣ���-T���,i�`$L�$�>�i��<3������ڴ�'S��H���>�P��*�k�)�k'O�ۿ�cTl�e���K���<7��Z��=q�2\;�����RI��.���%�t��5��z$t��s�����}�|
_�4{ծ�Že W�W��Mhш~�e^����E�jB��J7���% �@G'�1F7�Ys����7���?t�W�~������Q�jl�8	��FR�b�ЬP� u*���&1E��ou��X�
�.dâJ�^��0|����z�i	�+j�=���]OB�pڳ�,R���v��Q!Xm.b��9�B�)R��f����ES��Nlf��w��������/M �ͯ���^���e���T�ׄ�C���*���-9�⸪[3��	��t�+�j�Dg) �짉��BQp�����άWм 4�������$�+Q��-�p�XZl]�i��#�`��+��!���ˢ��H@�^���oy��ĽGl��l;�-+Ko,d51���$&���3u��*mq�����17��T���s|�a�0�:�� ��ZX�Iwu%�u����[n%��pⶈFȥ/������q�e��5��S ^}�"���͕z��,$7^�Q��ԕV�Z�"Ij��Ҏ����1�g@����ȓD�7��{�rZ��B�vF8~̋�P�� Gl��	���0�d�^.t\���q�" I��K=~<�DFJ�\8�TXlxVHYEB    fa00    1dc0��3$�^�����64��\�h`���J�U�($Ǌ�:E�����텲�|���цt�s�=\��'a�9J���E��,�0�d`H�5�d>^�|�@�~�\�̯�Vͺ��WlA���߹4�±,���`U�9i���S�,�
���h}�/����g��U�(:�I:e�'d\�p��&�;��d����S6c����� ����9<����M!�}�v!L��Q���r	� v]G���e��b�2��F����%B02���3Y�t��i}̀�J���ym ҿ��B���o��,�Ǎ�.**3rZ����j�pW�d�q

(�Lmn��(О2��9��;)]�DM�e�V���K�����r��\#���Dwj�Oᅟ=2V���J�_U�~V���?Y��|��́����=+�q��jwA�qs�K�mk_�T]��NR6O#ڵ;����vBXq�*/�Y�6)Kf�<�a���71ځ�Ikcr�-��rP2�7s��3l1���a�Vv���fLk\��˭�	
lm'�T�)/R*�j��i,9�zO���QSkiq<��D�D�ۜ^��7����K�mue]w^��8e�����b�&j拍9��|n����)SCM��CE[*�%�!��z�Uz��i��)Jsn�SJf�8�,��l��y*��L��r�7��(���U/^��.���Hv�΀޸��?[���u����"�u}�O��"g�d��)�{�2xc�Ă�����=%G7
s>v���Z�KD1����͘�������9L;�?@y���[�?nJ>O�u�Y�b`��G �`7X��\�ε��2�B�4��ل�I:�sl���-Y�����J"C�s`@o>p�<:� ��d�h1|n�ߪd-l�j-ԵzZ>\MKm�b��Q�%��|X9����ަ��k���>�Ƒb�O_��Xl�k��?e�&|����N���B��� :�[(���[�n�@�M>��<svJϋ�L<��5!�P�܉б����V����Y!�+Fg���FQ�79�?�43{�k��֩c�W��Ǹ��;X���8H�ZᄶHGH�Z_�1�?�Қ��bm�$��8���!���i���z���5y�*o�~烗��,0�!����@h�e�g��i�b�8�)�7�4փ�x�@�~hc��ǡ�g�=ؼb���1�.�3�1�V$�q�-%�嫦V��r�M�n~_蒈v�q�f���)^ہ�
C�чn�P �S����yV��z���Ѿ��1��_�������ft��l�f���}@�^��l1��O
G��@�-?�%k�jY>5|[�8���tf��X�,h�!�]�����0�;����CG�Du�о�[�h�Ɗ��0,(ͱ�g$@�S�c���Koԁ����]M�s�)��G�%ע_[�H���nT��
L�dF�#�qeT�^���X������p��o3��u���:�u�?|y�6��������D�?"FP"x
��c� �`�z����*B򕳏��X6�*��(�@��>��̍�- ������*� ��yoȨq0�W����D��m���\ĩ��)���o�@�(��M�n�kk��V�;���	v3����#^ދe���i��6pI��{�8dA6����,�=Q���#��K�P�)�}�~�^�ʳ���-J�f��NW{�t(}ooit�d$���?+G���V�Ÿ)�.����x#4�n�	����KʐđЮ��S!~[��D������!
�=�G�Fo1�
&���������N�_l����I�]�T�o��tO�0�5�* {r�[�M�2*) W�
!�к�G)�"�a� ��/8��v֐~'�u�2�]�Z"R�֋ST�)��#@��ٶ[��J(��\�5�A«i�ٳ�����k,M��r�}�mON�`����{�t}�x屘��
��Z��ƽ[x#���F%�CL�(�+���� �y-X_fU��N�|Oc|��^c�O!��������դ�DR}QQ"ե��!N5�>�U��QG�E� �u`QR%�ܳ�[x9QL�4�4����9[)l�,���z��Δ+�����%sO�Hk����}��L��;yx�o<y/�f�H�y�<��~׶3�^>Yl"F��lLh���S�筁��R�.B����kH7=����լ*J��2z���n�%r}�O�t�9Sﮡ�N`�[p�v]m����~2�A�i�H��T"{b��M�����sT���*m���܉���L-�X�z�-ĳ��ߌ����\��������]!C�����	�J��Td ���=E@�J�0�>hIN�N�ҟ)�-��d_�n��b�@>���!�^��_ Fz� er�@��o���)�h�2ĪT��c�����o�����+d�����_;ɬ`�;���#c��i�HB�}������8X'QlK,~:���;7��Z�0g�� H�� ~�{4��2[����@N8��	�;\]E�L����� u���$,�E��P	7���k�|�=;�B����ݛKքrc�|��j��|�ߝ�7��s������s��R��Q�L x&T�ݩ�'��	��I��i��cx?ٷva2���1\8Zb$���U�"��9m��۩����c��Z����\�uP&�1�wZH3���>��w�r=���^ϙ9\��|v�D�U��ԭ�ϰ/1�r�^0~�Z0�inE�⎼ū�<��a�G�7�<���NpӉ���h
M|<#Q���
G�`�땨��ˀ�-�];q�<p�o�x?�dW2{�����Y�{��������<%�P(+��E+W0�X�\�����\��i������(ӅP��K���2��إz%q�π�-y�)~�?L�9r�F^���'y�ۉ���^^�!��@#�U��hY.3`0+���2~V93��>dˬ�Bv qL�v����6���<���$�j0I5��$Yj���-(1�k��N��Ԇ��}�6�Ϝ�g�|Տ��"�)|��w	~�k9��´�%�C��U�h6����)�>:�x�ZvqšC!y8����6�'e0�<G3�(8���F���6>��dEkD(�)>Twa{1Q)'��I�H���:N2���M�%[�V�CE�X��ܔ�~�K3�|K��d\7|f������!�A��(��D2�8�D_���S$�a�>��IH�!�����E5Bt�ˣ!rj$��M�`H�C���Di�
��nkGV����>K.M�9F������3��5����'R��Ѕ�$�d/���Ӏ�ߎa��9��S�8}���ܱI��We��F��u�i�<։��o%z��JR� �b-�K,h{T��LjV����a��R���(3�E�X�n�jʴ>1�G\������jY�§��b�J��{�����Г;���2O�S��*;�N5RZy����C�+��=���JR�_����H���ǕZ	R����KFg]�*y�R������zU��<�6�+b��(������6�t� O�D�x=����t���i\J�נ�hI��uLo�|)h�&:ȉ!�T+�;��0Xb��%��t�����uc�j
�oC�d��U�����	_�J�\W�"H����q���"9�έ��n9�5�3��ۮb����lȋj\I+�m�ZhG�.GY(ڻ�Q��0��nǣPu`����,|��`#�G���C��5P�����!������*�*UD�a�Ŝ��B��%��n?;��vk����P2=iq�=�`��߽.�T��O�Y���(�V����ʉ���B�E�O�z�(h���������O�F�F�_k�9���l�M<���X������Ӿ�>�Au�#���iځ>d-{��!6,?6�� N���zB�	�b]q��#'+3Ag�*V5%ǳ8���Q��m��d��8��W&j1�V�xe޲-�|2�x�+x������ݔ�N��S��n`f��)����,�n�����5b"�'�ԕK���~�"�z!����+P�qb�0+ 1R�y3��C'� j�Ga��حm�y��<�#$	�e M����5�myZ]��Xp��y�'��b�@���o���a�"4Xz�\��L��Ӓ� z����+�ǂ�ͱh>�4t�ڐ8���^HډT�SE��7��#��c<чq	ywMk.<C`i���>F
H�ԴN�a�����3���,�G�x��~X\L����u�н��%���X�8���{'�|�B2��,�R;��a�DN���O����N�Ĵ���1�L�����J2�0��p$�n �<ds2�Uͨo��������P��S��������<�����ՄyP�)]j���ڄ����w��y~J��\�|�p��J��)�Y�^$T�ֆ���ؚ���z�����du�V5D���4ib*���-�pU��\%y�(��i29�Í�m)�"��r5@C''�'i���}uL�"�>�+:���*�q���@�M{�K)��ȑ}?1��"!���S��V���D�k F]������7a"��2n�i�jA)�a2���fwB&@e��_q)⹳�7���na���<6��,⟎�Cg��T��I�J������YICS��.}�1N핑�0��g�4^R�ZuA��ֻ:���-R�OS̰��s�ך3e����0p����=s�u=Gi��������ۭɓ1�.��s/ �Bֿ�F�)�<.��v���$��J�Y���V�����彴/,�$g[*'�w�RSL��Lߢ~]�Fc���ي!�4
��a��[7j"5��������j�\�T*�vY�¸���v����C��|�,��ō�d*v�{K�Z�n+ñ:V-u�>dXf�b�YU%�NP-���O6 @��E�vw��#���G�\��Մ=�x��:�'xp))������5��*���s(fp }H��MuJm���lb�ԃ��3�mHM���V�S�1�h`E*��&��G�6t��D؍�$�|o��`��pz�y����F����n�qq�M�J�=
3��G�ǰ�2�g�B�u�X�C��p\���-a��iBp�{�d�+���(�/�V�&��"9$��4/'��C�$�'O��V�Q>)P����GשMT>_�^`�ѣ��Æa��ns�j�kg'��pƎ���*|8eyh�	9�J���_�� ��oKk#���u��ev����}��Y���zI}����Ւm\�̇��hz���'�����q��b�C�Ty��"�����a�g�Y��Q �]q�eKA��ɪk��t��q���f=ٙ7ˠ�t��J�ۋ��`�_��wr˞Tך!�~���1�O��PS�m�O߀o 0�����siY٢IoA��:�Xb�ao������M?�{QM��U~��b��/�n\�\\��9 3|�,���fgn*L �7aYee:�G�l�X��}�r��K۱�B�Ͼ{��f�^fz��~�<�./��r!0�D�z�p��tsM��d8��X�u��g��~}u5N���Gv�<�c$���C��9����8ꑖ#�� $���[���a�3�l��u�����č0ȧ#!�[!�������7y!0q��߁`��w��e_MJWC[��i8F�:�U���H��k�7ӟ��ޥ)����	�����Qz���d�K]rO��*�C���[�t��j Ha��YP}�������P����$��;�y���TOܰ��cX���0,��қ$��bd;'nӷJ�.���[3��O:>�cϖ�E��1���u�N�u/���~4��#]hq��`M��6i}UB�0�%*�@7S���j��8/`��]��w�{�������n�H�ӳ�I�Y����kG8��{�����qF/t���������yv��j+��N�>G���mW��/���r���6��;D ���jY�L5����U�:��`��ѹ3��k���GW�nx�3gh�ջSf��Qa��I�RRL�����֘L�6�����\�.��nl5&�~h �4퇈��$�>�����j�j�Y�>e�/�?x�n�O}yv���F]eF�Y6�_�שj`�\y�,]�>���0Dl�,*�>�\;~�G��x�0�T$��Whƃ�����krI���B9]}���苞�ٽG	��!F�#V�K�74|9�ܘX�.�<8���4� �B([V�JT�M�g����X>J>�zp%BPq�{z�#�qj��&��e��# ND�õ�B�^D���I��
@|iq�[G�ǖ��=�>W�ZEҶ,u��ەЕ�8�!��M_Ɓ�C���_΄%yۭ�KW��>�T���i𘗕�L$Y��P}�JD]j��@Jy��2WXuK�i������C�{�m�2��s̬ݴU���Q����_*�Z�J;r�L�hĺ��HA��Ї&�����8�f-ֿX���<c�����ǎ0�12��,�;z�&���r͖*��f��e�ЅΜtf��)��\�u̢�8�\�ʋ��d\.2;������fnha`�����>~l��~@ͷ��/xX�,l���f4�<@���æ ���ʼ�M���zi��o�P��C�S}����s��O6'���ˋ���:F����������u�ce4��������y9$ަm�a
�$��#QL$F�J���鮛�Ai}��y� ��1G�l�;�L��e/����9�{�������̕!׉0g���]��ep�0��\�T��;�/�)��԰pkPy�ͧ���g^!X��`�T��a����Ut�?G�X���{ȶ�&��8T���:�j�4�7�ֳ�U�\%�2��7oI7�פxu���%�o���Rm#h�O.��b�c���^G�v�ѴD������`m+�A�:T!~�֭s�!sVG2@�Y�����ys��DˊRD�$��0�.`�E�@�͊!6ȕ�\C�.�F��PN|z��~�3&|���]A�<8Wy��qd�����Y�=AlE�l�8�!�Kk��G�9���p��@��(����r�>����|��&k׋A�c~Bo�0�g��� Pǻ���Jc�S2q��m7�/�N_�⿹}�������6�Ϛ|[}�6��\�"6�ѹBj[Uʹ�g�H!��О응���9�څ>wx�Xa2G���"�[S��m��3�ll/�xFB�VB7@x�����W`ׁ�!�b��c�1%i����aF�B�8��3���`i�#,�E��>[X��m��/���5T��zdb>�����b�țND9ϑ_�18�y%>@���(���U!ɝ�Lv�?�pE53��W`5�[0����]��5��WU�i��O<j��n��9��U,1L�u�Wg�;R�Ǝ�C�_���_���q�\ExY��[�n�%�N�2�=��p,�gCE$l��v�XlxVHYEB    e7be     d80�����|�)��p�b���j��	Daf��Uƪ	�fa��,���|Lv�f ���wZ�e<���酶zS�q7,��%��p��=�i�u��@J5�^��}lYmR��sümϫ�"�[S+D"{99{�� Ŧk�r�.t# ǽ�ё��e�$x�]� �an���/�]7h: ���"9l��di:�͏I�+���
�z��HӫSְlƍy��`O�s0_�كO��3��c��&��Z����P��V�f�2f�R�Y՘QXΏ,zR�3��|w��g�����"����Z���=���
y>z��@`*q��h��ţ+E�G>�ap��֒&��5;d' ;���O���iq�׎}�j��ϞE#��^[��%��
wx�~m�<$�C*��M��7�J"�W��S�HA�֞Z��Tc'X��������F�6᥾	]-O����O���ٙ���߭US-�F��ę�U�%�X�.�]6�U�(��1��;T/�G2�ͬ{�o�QB�jϠ���bO�|F\�5z�v�̘]�褓A
��tN����Ǵ����al���H�҂-`���6�R�5ێ7F2m�B�H^���h�/q[�M:	=��Gҍnlr��}����u����h4�m�hy�7�?-���3�:nUP��ܭ~0��c�drk��Zv%۵>��a��@Zm�^;a�ń�1i����,��P�)N?�K�nC/�2i�n2���^���t��:E������Z�KȖ[9�j�к�މ^�H�a+��s`m䏯/x4���P?������� �9<�b�R������Nm'��3Wӳ�~5m�iLhuȍ�B��4"�Ja�3���f�E�bf+�qu`5@)���1�v��]b�I�W�����8*�)Ym�nF��}�E,�qn��xsV����^�"-ˡT�
�}�!S�+CwQ��!�z�\prP�ݍ�F@����V��N�$����͇R���VB����5��������d����������H=eD�Xm��+2a\�/ M�����m�!���]��E$�nO�,B+�'o7P#��%�eu�ZRL�u�J�n~D�W���W��N��� �y8�Ly3��fZ�� *s܉0$��Ƿ�\���<ezF~��=���	��T$�!KyA�, �K�h~���]#r�&�X5��ò�K�ϳҨ�!�t��C !*}�F�G/�=./���4����`Z��N���i!��s߼��*��czZ�"U�r�*��sֽ�3�����`?��x��_oh����{ר����h�ו!x�r墀�nd�������yi+�c[\�Q@���R�x��V׺��4�|j�� �\Wd�{�T<�1.��75ah�-��daz��V��f��ҝ]w�N�Q��A����@�J�Qwl��$�l~����[���}5�&�\���ῧU�?r�9�� oH��I���� ���3�*�~��P�s��bI���B2�b�B�$)�g�?��0y_�ber�E�L�s2�^�y��&i�-nH+�k t��_���$og]���M�eh���B�
{����²I�C��;�g5ٵDL�8�~�r����iF6.��W�(�9͡�O�EB��Y	��0k�t�0Ү��kU1OD�$B�Xpڃ���?����4E`��ű�"oIh��wN�	(�����}~�h|����7�I��?�����R5�Q�+,�T�H�g�g�3(Qj��J�����Q$�����N}/��\2��ȇ��?+7r�A�"��� ���6�.B�J��w�2�6�V���=�ڷ49&�WbġU�h@��'��x���SQbX�3�v������
�\���듀耘�\�}F���7{bֈ�+����r�P���$o�xn�m�Hqx��O�a[H�|$(Ӡ2�>�ѣ����a��@�14�s+>�\6~�_�|}gʨDzk����J/Y+������i�Z�l��W��T�Ì-ml���>�����åH7�}w"���'9ߌ=$ȇn��h�	���ۿ�����Զ8�le�>�˜FB������'�� 9�B�rW �Bc��~gL�D��e�c��.ph;��$�GQZ6yb��������f)�/4�cG2�С���n�a9QԷ���������{��U��9nd&�b�ˉ�YT/U����^Xr�[�X:��t�a��,���c҈�D@�0��8�ۏi�۫b'�r�j7�~I�|Uُ�lF�"i��P�&��JDC>�� gv�bA�˥��}�ˁov7��_gga�����$��R�i�rM|����7���L�~��������FȀ)y�nDD�r���e���!���6�*ᲸT�;�S��A��u�F�����a��i�e�����p@� ���A��)��,��R��\$�|�d�;���J�%k-Ԫ����_]���
�������C�]��z��[I�2�+��g���m�h���YΎ�������I�!I頻5zt����Gf�_%ፈ^t�Pk�]��s�#�}��ݷ��kS}�I����Si�]�����"�@P/�R�Љ�("L�<�Bg�^ �9O|ZȌ�9<z͑j�0]Q���{;l�`T$�fY@���0���k�^��K��$'�i�[ey���D9!'�vt����~D�O���J8�����h n�b=*Ȱ� r��L*�E����Մrq����<�2#���u#�x�<�t�?���L��ጽ�䴐l0k"0�����i�?��}~#(���v�$%jG B�'�M��\To���Lh�U����	���u'u�W�2"n�z��W)��4���
G�Wv�eNپ��'(}Z��P�#�$󀻳Mc���do��>�,��f�Rբ���'j�bi(�Ł�+%�~��j� M���=2�}$�����)V=�zU!~�{w�z��-{x\YR��x&\oUnOS~]�)n�G��v�y��Q�����&�z�� <H�6y����|�K�X_��mh r�Q��i�7�D>�Q���\%ô�z�H�ʏI��~�v+�#[4��Y!.=�T��h�4���'̞�AӺ�BP��'�si`�������7���[�p�i��<}�t+����Xk`=��ͦ3���}З�K>ڞ�)&��
�ZO��!eN�c5�R�~@L�e�5�3�n��eR�j���[FY޹2�F���FRwj�[ݩr6�*W�kK�cG���F���^��(���]�;�������8M��_ ��|PQ6Lj1/:(KP�ʬ㐪M�VUxjr'�܄������N��k?�2UHZ3�,���B��D2��O����;X��|��!��po��(����ͥ�����Q�c�7��"I�`�y�I��x��Y�㥇���X�0�E:;KG���%Q