XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%9)�즚�7���IL�P�ǵQ��TVH��]��nZ�Dd�*nj���q�I�O]�������iL��C�^�,��R;@3�3��d�#� ��^W��1�2.�8��h@'B��`���ZA����C��SN�u��_~�+@�k�iܜ �&~d���'b��+���+;N_��33PqU����S��v�'��'�3���֢�|m?��u�=!�9�/;1�)I�ܼ`�3��~��H���<f9�������ȇ�l����t<��+A�v�j����5����|��X0-L�����sH"��:3~ v���nN%b�{�%�U�3I��s_Mm����)URT�zL�{ZvȚ%�c��?��LW#@Ü�茺��|������tOXqI#���>ڋǫ��j��xL��@��(�x�u�yԙH��حa��?�'�ߪT�Wǆ��m�;�2� '�L��!�?�}�hͦx/i�Z%�%X�����7���Q������`��(1E?��M_%TF"�wO�.�vs�������=tw�R��d�i�j�����jJ�1GY
���$i�_���$��a��%8�#c�p���"�p���e�6��G���6�1�8s�A��@��*7����G�Z��#sH�n��@ ��jλ\3�(�_
�l�	K��%eC �F��&�)6_q X'8�1�38EN׾ +����)��~���W޼�P��%�5d����%C8����U��5��G�:�E�� @�XlxVHYEB    dd8f    2160�$7F���p{�����Q���M��_��E��7BaS�|�Ш�_�J��c/�ۭ?��̷b1���	�Ť1q]�����+]��A��
�lL7\�c�@��$�S���Q��P�;�ٿ+�L����E�� �K�7����,m����4kdna�1LX9螛�=�aB�Z���N�N�4)�<GÔ`UM���o�,��!&!4����o}|F��In��?T��.�x�~�xdjIV웍2joa������H"T�{C@r����Ų�����WMUK�x�����	6��5A��d�4���LKP.����a0�2`¥)3�W� FGD��s�߅�%��)��]ˎ�"-8��`Xh���P�=v�V���]V�2�༦�x�|�6�y�|����d����8+%�(B����IGlE������-;C� �!�����Ovb��L��p(���m��Ge��٣����0���z�-"jJ�x��z[�1�_c�]��Z|�d��L.,��t���&������i����G��2��)�-��o>҉�JC-�F���M6k`;�+`
����X�=�I	I�u��W �5��n>�Ch(�IWVa���Č��\��y�N>�юe��}��r��Z�΄p�߉cD�� �_�jN��>��=ȑ��u(cA�5�e��v)����|��yC��ȷh%�����_l�<㮯	5?�U*yi,N9�r������R��W���N��=�^�$�S]������e@s����j�Q˥����m^�1��{2�<�ђt��cA(E���c�74���y��%V��\w`�ħtJ+��84d9��e<�bTHtgnoA���	w,���[������GW���I�oM���s�@�� Qӽc]iM���>
d��I{(���栮<!w��@��W���jLXND�Pۏ_c:;��:vHS=���Ms��z�	֙
:��1�1c�aEH�A��7s���O�/��m�_"���3�Vl�Qx�2yd>P�c���`��z��.�:��s��1#/�4G���y{���Қ���<����R�Vw+
M�:4[����>A�8P.H�-����_�ΑD;��@t�5�����7t�:J��G@�I�f���ɐ��{�l��'${.{y*I|Q���r��Z9�rp�b�;�X��=�j�%���1N��~]V��^�̛T��3�m�ގ��r���9�>��(�F�(�ja�t< �e�rD-{�;bRY���_29��rU��kL�q���Z���0����y�S�G���A��g>:d���G�������wZ~��ZG�bH�'�Ek�@�PDJ����n ���HSq�VG��À�UN�����0�1�7jg�������p�m
M�:M��f�I�<�7+]�L�p�w^�?�]��\$�x���W+��>q	S^t)�y�5P��5S��]���tL��V50ś�E~�D
�H�J����cP}O�$�MU���Ǯ�/ڣIu�6���ɛ-�P��z-��Z�'�C����غ;�� ��u3��6�V����F.��K�
�������ݬx�j7�U�+�W�Ш=��~�6�2�N/dnT�zq��`�@�|�9����l<6��˂�Y�<W�!dWU�Ϻu�i����Cd�&X�Va����J�Z�"֬?��C��m���Ry{��4:EIV�M�?��?x=.g�~��DU�瀜��;�3Z�}Y f�K��u�+�Q���ϝN��$�y�W��z�g=Hy��E�uB�Xbz��ՙ榏��z�\��=�]�#q��D�GG�gi߱���Gb#�l��Vn1�!�Mn�Z�H��)m����w�2���-�����$�����r��V�[<wԘ��O�Q���L�Z?��.:[X��L�0�8wc���tl���t��֏T&n�{|�;I�I���R�x���xC��SI�\�i�Q�����`�d�5!D#�i�Q�I&I�����������-I{����:bu�e��C�Bjs�]���i�n9��h��&�$t_����� AI|����s��D�#%/�=?��}Zp�U�Ր���=d�C��:
�'�ה/�ToO��Z��ͺ����qUro0��{z'�Rޏ��u�`���f,)���H�WOAhg��<eI�Ljx�e���nL�ێ˯k��ׁ!%S��u�H���!�x�J�~?׃n�_`KY}�+ʞ 9)AV�8b��G�w��(ip�S�+�������4N7���٣�m��7��^��ʙ�0]���h�p�<��m:Y��8#�G��
�A��ڄKk���"uJ���@^*������&�����m��g���/�!�O�Y�(�얰a��GK��YFc��`�u�d����~��������ffE�w�y��U~��{-�뢦i�!?��ð�A�YWant�Pk����<��x�f�m�)K�_��F:�Lk'!k��M�ߕ�o��-(����������p�y�!,�@.�u�9�L ���.L��N�Ո�:���%�A>�<V[&Y��9�P��Eڗ6D���t��g�X�'�J :޺�{e�R}k��pbo}2�ݘ][�I6�3��Y�y�܅̿6x!�� %��p�,���^���)��R1�����g*��vBY�.ˈ�6��B`GGYz5�8K�����w�@�/��cG����DV��;HF�DX^�h��rj;}'̮WoiL��N��SX4�3V��2ˈ�T�T�q���9�{'��5Hj�d�M���ݳǖ��X���[������3]�ơ��Yl/�������v��Oq?����<.�j������|Be4DM��3	�Z�~���n�����e�,s �nLP�]eEҶm�<<�o��wrH<�٢��N鐐�K�>kYA�|��^�NE���[I������]d�Ǵ_�����a:��O%��<�1z �`Z({��@o��wߩ�6��Ј�-�_�WҰ �(2����H|�eS&撒:���ѶXx��)S"P����K��㞠��d��x���VWb��.���ג�c�����m	���b�`�b������s�|�76;ƽ�_��%]G��Mu�9�����E�ؑ�	Vi���Z~ը����U&3L61����m���>kUVc��xI��"1ϡ6{�;d��@��)@l��s�k	H�i�'mӗ^;hK�0�<�<I`K�7�Y�Ӽ(�L�m}��/9��?��C[�o����$|�Oܲ����/onr2 �+9���k���҇���o�_�2V��|�#��/�O=�ӝ.��(�j�a���a�V���3���"���8V(_���ز#S�������tۛS�\.%�j�5�*��ÚOη9�X������#9p�}�������GΒ+�����n8�C���]C��k��x�Ta���eN�O� x��@)o.��-���h]|�5ք��kN��^Up����S���cψ�դ!��M�����`����5�u���=nE�D�����z���S�S�]�U����*��C�"�|�j�ѐ[�C�e团9{�p��҅��'e͕6p��i�v�2���H���1���M�;_��,�縆���K��"��Ni�����X����I�mݦ��6��kЁ�FzU;��#�HrE͞~��Gɫ�Vz���;�C�A>E������bnlcT�Ӄ"�a��o�vꛢ��������58v-vJ_Zs)Δ^Bw��������\�	hh3|�S/Q=�}T$Q9�b�fes�}u@�����q9�0�8�4�&��\���J�-�Gjj�����ڨp�ԧ��,/z�/�^�}���ih|�Q7�)̚A�;�A_��B80$,�J2����X'_v{�\�(DC����9u��e�8,5�o����[uX'��dJۜ��Bb���3�E�s��f,MȌr�JWp��兩8A�p��l���d��oi>=�| ��Y~1�g�ʖ�0��*���W��:�d��������Vn�b�DX%r�Ŏ�0>/e�䐦�������"mu�/���������m[�o(�����'Z��n+���P�A��O���ZX�����O��,o����5(��kzc���Ҽ�i�<�#��hb�V��4�^1͋�������|7�yք�#L5$j����cŏᘿ5)��p�J�g�&J���T�0C����
�~����o)���_�E�D�A�tsF��꧃�`-F�.eǃSԻUhB�V�n�3gV]�O����k���m��eG/;�:�v��=\�@�IvIp'shm
��,r�u�����"�v���ξu�~��|�����f�]n��2��[�d7Ԥq3�	F��-5�)�{X0*�&���W{a���Џ�#�g�#g����O�ۙ}��j(j���@Sц�1;ԑΑ�aݲ��Z�`	n���GnM���a��&<#�d\9�g�)4��/ރ5DdG2!ߢ����&�Y[�v�_��/�Jƻ���rCW�5MG��/I�g���^����;��*v�Ũ�������������y/��Rl��O�]}f6�D ��r����;:UЛ��E���1��t_��Q}����c2���U5Ւ������	��+�}���%S0z�{������^4�G�c�`f��3ӈf\7�DzD@w�8�y|�=\/}{�	k�9CAt��.��]�D��8i+z1v��β���Z�@��閞X����UBeD�y���E�N5��� 2��h�fRS��6jUDsJ���:S�B�_2_v®W>�7�����H�!c����@ܯbYzԒ�ah�>_N��#�I�|�2���:�O�V�\��5ؑ�X��@�s�%�k��[����O�3Ŗ41UA�T���f�X*���2�2����&��64"}��� Gl���B����e�{������$���P�6�9mh��ǌT��A�a��G�I���X�='16ņm�3��`��_}$>����� ��*��?.v��L�j�,,�ڭ�O�/+}���a��� �� .>:�;�=��B�¡޶�S�e�g9��Y%��z���`�������
N['���W
�lck4/����!�y��#��GRP8�5���4,d��e��M�{��rp#� ½����
�KƍU��V�s�Į��J�3#Pб^?�E����H���������B(��7������/�7>1��(`{��U� �b)���k���$��A�ӓ��_�_>�3n��ۉ����t��h�w=�\�U.�6���M����%R��X�0f�:CS�n��M���#�/X�����9����5���@Cb��ar����iW���V��HՔR���v���"�q�tMp����U�	�U��Pv��65n�da���k(�;,�h�{��W�[��+���ξ�GɚB�{��:g�mq�h�_�=�O~�9'	�쾟��|2���������*�� ��A�*�<��)O��L��[�R�:�Ԭ5
��ӌ�W����18��qX����|���������{�ˑ�/lG��x�Ӓ��Y��=���s���(�7@\Y�q�n���Y<\ ؍K��6oK�C,4Im3\Ă>�S	��!� �w�"B�+�"ρ�89�$t���^ޒ l�Xõ��
�'=��v?�ͅ�J��������mM�s{�}�94���������k�0?������E�l℀��	z�E%�xM��}�F�R�@&�WW�dR#�C#MP����	�ѨF<#��R�8�]Z>�����rh2���>}:��,N�����V*08x��E���D��.���߷\�j�/��:�/H�3a�����1'�˱�����ʱ!��-��\Y�д�;��Nx�Y��};}�qg^F�l�ռt��gɨbo�(U1�^��
Ч�ȺzK	aǬ���п+���}�`.�x�ݥv!ⱷ�KnL[��������V�tXUߚ�޼�k\lsEa	�)�mGCq�fh��HU�t�:���d�w�*�����*h}���rp��˫V#�uI �H��LÏi��3�Ȕ��$��-������\	��R��{���OSg���mc�t+�ѳ�NP�x�����QGU�D�B�ҹ�]�|�q��G�����e�9Ȱ�ˉ�m�,����)�!Վ?�����Ɣd��g�N��< %��J�0��ޫ�c�Y(�Y�2��6M%��R�T1�-�bgvL������A��0�=zAO��
�eY`�<��@�wI�9A`�k����w���Y�r��Y��^�p@S��{�=gI����1b�H����{_�RYa�
"���4�����O,����X�9���}0���Hp�}����aҼ���ya�Jg�'IGeX���?@�Q�h_�b�?@�/oJ~|�V�wޝz<�+�n���K1��Xwz�@�bkmtG���G^��ݕ���Ѻ��☉�w�W$�T LT&K�H���]�:� l��тk���=��.c��Rx���08�z�/.�5�I���a�G	I�%��0�GW59���IҾ��i�\+Ժ_Tp���bgi�Lg�����q"_s6ty���F̄{8݇���*���d�����Р��%CQ�
���0l3V����P�_�8mfJ8�+��##;�'�)L\|�������1�X�d���/ Ok�O�YC��_�ZF�<_�~J�k^/�%[k}��_[��Xݗ`�d��d�k(��\�|��Pr{�z��Z���Ƹ��I�:�,!W��8�3U�;�������gYlq6���_]_��f�й�`��T�3�Zx`�Q���� �S:�_!®/�^�x��ʤ�����Bmsn����pN�b:�?�O�9��㵂��?��%�I�q��R�D��|^�ݲ����o�(9�B�?����Y��A��m�t܎��ss�װ�t8ܤ5�U�Q��Pl̦F���\�B̿q��"��]�+G∭�HoOA�P� {r�Z��;"�@}C���O�@�UL���0%�����l�^~��c�KH��Y��J�W�*����a�j�WپXRȜN�ѱ����_r��m�Aw񳸽�{07t�(�3e�a'G�*�Vp�����PD��%�����*m�"�Ϛ�+��|b���b���Ҥ�+��	� ����`��ʁ����1-u�����O3`��MT[��.>�����>�G3
Ρ�ܪ�lL��:��8a�*WkK��;�G���/g5)V|RM��
r�\~�$ƀ@�U�'$��U�"�Қ���y�>�ϹgͳF�κĬ���~񏂸�5[����1[��@���h�?
��	�ڵ�C��zY?���ݍ�o&�lO�P�E��ͳf�v`�/\5f*����4�)D����"Α��\}zA>= �����r"
��?��dv��.��u��dl}u:���{p%�H��w�*{Ƃ���Z�����R��Z�0P)=�<��b�WJ�a��!���8�"H?���G��8ɠh<��6�c1��'3NtR�����7B�D�yshҵm���%�d2,Z��1nR�,�a��a����%i�`���`M2�.j'���H��2�dA�&2X3��Ǭ�,�����_�g��_H�p5H�z<}�8AY��$3����vG!~�/LHؚ���Q�'�3M����ɩ��Qb;U��ՕΦ�N��Q��(W�MNW.݃��V�ɽR:�v$�i������0*�lY����ox��CI=�K$��`a���� �=�-$F��I�e��I�U�o����e�ϹBM�x��CC'�*K_��&_���8g���J�BFӄ�f?ٛ- c�e_%e�C���[��.z坏?�L)�X&��y�@ւL�Hx��� �%]	����PpA����t��7'�AR���Z��r�E�ӡo�����H&�~��	w���2E���1n|K�h���m�i�R����'�CoU����!��[&������P���0Ӹ�lY����y��"۬���d$<�nvm����Ҭ�^�sVjr�n�rz(p��2jP,��u]�L5g�}I��鮣��k�9I1%L���<�Wċ�f^�ß?�ytG�(SQ���)�K{�������̧���sD�_���5s���t�&<*�W���{+�<v�F-���A�� e���e0�K���'���t��|��br�fh�ϒl$��*4ҡօ�d�<"4�����J�˔�@Z�:]i�J<eԷ��z�� КI�U0�T�V�v�I���Ef;ˆ�~�
���ZˎC�:(�