XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|�km�T����t
�F����m��i�_^n�ks�n��>Y�Qx�~��oKɭUjY�f0>˱b�Q���`���?CzU+j�m�^�X�)@�o�vy*�OWb�j��%�
�K��uy���M�j���R��K^������@y��ߎ�����'�o���J5�P\��(�X���N�m�����>3r1�J"�rS��)��,*HF_9G��j��uc:r��Zo�|$gP����&�Ҽ�$������/&\�UIQ���+��aEAU"����?+����u[�Q��R4b�l��ykw�ߖ��p�����%#|�,��}piqV���㗪�����6��Ǽ[5�֨T:있����\윞���j轴�`HM�x�x{��2��S�í�Y^�F��!��_r���}(�d*��R���
�Qh��P�dt�Qa��b^�Oh�[�§��c!�d�sIcmJ�Rb/�A��ܓ�T	�!�F�d�l����y�J⻙s��-x����(-��|�[�K�9Egdʐӯ�*R9}I��A���������^����^.��V���?a���x���u��ѯݟ_�72船sfͯ�ⷭm����j����(di\���<���&�~���9"��MfT4/� pc}΃��a����31�)ml}&�~H�W�)��p��w�����U�$Ԥ]dq�\/>�(F�O�g'��(�B����$]i�Ԙ�,>��0Ժ�������C�d��<���eQ�"�qZ��5S�y�<�
S����>XlxVHYEB    fa00    1f10�r
W^�^��Doca�QQ����Y��NG@��7�P�]��ٗ��$��
%_���b��~ǱA7&����Xz�T���j��_c��5���)����(i�mG�z;���s�Qx��-Y���Ä
�zb�A�ٜ��ӈ�Ʋx碵� ^���H���$S��L���,a\�菺�&��݌_MjΧ�UL�!��x,���\H�8��Rb�ٕ:�]*���^�*B��j�n��n
��=c�� 4E�hpZ-��UW��g+��I��������!Io'�	i���ja����fM@}S�6.R��V:����/���]MH���T=��sΦCa|���чߖS�l	m���-CO9�����ю�J�e}�鴔,n�3�&ë�dN�<H�[v�މ/LB�'葇fi��;�����w�IX�@ۨf�{V��F"���`�w�bs�3ڣ������&�M�?�#~�M�.K]�s�Ԉ���8%���=<d{](m���n1�n�D�ѐ�<q�k[xY�+S�Ʉ���^�J�E � eNx.���+/�G.=l��3Z�_U��yq���5��z;�b��x�H6i�'�%���B���17���,�� =��7�L�RR�2]�7GWr�� �#aA�_ˁ1b� �MK�A�\�����
[�l^1,���=9 Z��F:}m�l�k���E�;b�=%�ky0%*S��d5���Z�C
���Y{U��Q���I\n��e�n��b5�~�KL��Až�G��X)_ӂ7T�t%���ca�ء%������I�$�*I�A���L��Q"�߄��]��O��� ��L�_U�&���c�U&��]ǒ�_'2�$�A���p��p�Z��'�%H��$�cg_;�؁���8��uŝT�P��	��%R�z_�oL�g�:�l-5�]��� �Ѷ�]j�uf�,9�>w�{k�Yͣ^xh�G��>���n~���½C���S�_U6�[�B���l�9�<(h{$F�k"qX8���Gw�G�����Mk��(�l%~3������s�4�;OrM��b夼Q(����W��	� *F�2nXKh�d����)B�x�{�&��
����-�ݘ��dl}xUm�3<'��Ɖ��!]�Q�3F�p����N�'��:[ļ�6�Գ������yP(3`�6�2Z�O``a���i��/��nm�bP��(�?U�*�0�4op��=�����s�i�d���;:��
�~���)�l`�]�#�O�wa7gW�/1d�U�gX�Y�C��N7�0)�j �J=Y]&�29(����]1;�A?��Wℷ
�{N�U�M0%A^s��&*�<�Ի/+�/��i�t���l��8\<�	FQ�c��u=E�G�����'Z4��n��l���Bii��,�[KZ�r٪����Z���iH�aB�r�N�f1Ĩ��#��E��J���ƺ�m�^���P��kp����mQ��B;�V���띞t3���uT�!ݷ��9�[�+PID~|�M+؛��������BaT8�h�	��=m�jI���lXy�`�/W�b� ��}Z���C��
�+�ȏ�Aq�(l"��i���N���mP��m]���}?Us���5��Ģ"�b�G�x��RS[�7����	i��طT�f��K59Bf$%���g����d����V�����a����f�V�g���M�h��r^�\�=�|����f�}f��E}EtY�Yx]�v�Q?j����2sU�e��O-N1N���S2�J�h��k��g}ڈ`Y��nR(U`.��B|���Cq�u����������4J�8�#6q�[V�=��Sb���q4΃�GL`l,�q6"���<����q�%~��tpY'5_ޟZ����@p�硴m��lw�ֲelb�sZ3�gR�D=��`%��{�:���7$b�=H+����H�m*dE��V�p�]�K���
�4dcƷ��n�"?�+�R�Fa�:�׽�В�;���u*w�2T�1�4�Qe'1�M���vʙ�g-eP�HXs���+S �=��M�қ+�+Q��h:g��Ρ��˽FI
�P��g9m���3eHe�5�FI\���g3�S�U�s��>t���^�Ǔ����H��v��K�9�UB>NO�@�����v������̉Q_
?҄`#�g~������vʊ���3M 8p�Lk� ���6L�
�֧4:cW��A)m�j��lA��r'm��o&)&��9�0U�F6�� ���W�:y��= ]�#�^����\mD��^�⇋�R��#+�ȷ"k�ks��F\�����h���<�w�5
�()$��red5Ym H�֌�l;`0u�2#�����r3-�d_�y�ȴ�lϋ��e�-T�y��*���&c��,,��x<��zHV�S�����!�Q]_
�����T�>;Ί�&0�K�lG��U�|!��E����ymUx��G ��n��(����E���u�� d$x)�l��`��@���[�ۘ܏<��AX�Q*��dZv��"���řa�P�r�7�l/f�>�k
~��|"��c�W�?|�Q�9��̦��%���3�6��9����ߟ���I��eܴ'M�1NqП�ڪ��l/nxxc6��E�f�|9A8_`�>Ϲ �y{��{���2I�d���z�u�]AP�_w�-#������\��̬wԱ8�T,��4�3Ĵ�R�F�gr�̕P ��`?�W����ꇪP��q��.�����%�S���N"
������>g+~�����|A�]::�g�8���MИ����>t�PY�2� Q� �NF��-!�GZIv4�9�� ��r�|�fm[r�ɵ�0�"�2w�%��2�g>y���wM�3���U�XXu��r�M��rO��=������'�"%���%�m�m�e,�Q�O,����3;,J��ɨw\}���Pd7Ș���?��I`*㸸=�]&�`�	�K��.�f#����f��H�F8Ir1���~�n/�u�l��4��!�\�(����\(��4��c�4}sU��gy�
P~�9 �CV8[^��v��M�_!ޱ2;��S��"5��˦��e�U{���Rf9[W�3k�!�hf����M���8;������{����=���q?$YƔ���E6Z9V��By
4������ÚSʏ�+�E>�[x�s|3ʴ��_�b*��w؄��iΣaV�=���n?�5���R;�q�����ۊ���\�Q��U
g{6�HB {��� �ʘ��?#D���X(�i	����bArkA1U����ϖS�k��9*<R�O��V�r0#���B���{X4l�J��v;���{i��,y'�[��A}(�"�H0���)ٳ�Iؼ�S*�&�52�ժd��ϲ�.^'=�W��d��!d����B�#\��b��^kGϨ�2]�f\S�?:^�hn ����4j�
�p.����s?X!jQz��@I�q���&�+�%}�*��2w��O���x����Q�NV���˅/���%�Q><F�p)B_1���Z4"
x�w��"� D���5����5v��x(��?>֥GA��,�R�s�m�~���@ߑ��u &���nV~[m
�%��O�R+��(����5�0I�eA牅�8��v�W� �z�P�(\�CkNv����K�y�}�m�D-8b�OͲT�k�� �eo=�>	3#^�y��!O�64^b�r�r+�%���1��_>��+���z?I��đ��c�7K	ft��YG����ĵ�.YmZ�h8�d:�z�p�~�F����"��y���[	1�y+�Z.����.����h!����i�0K���|k���� ����8��X��LEt�����{����%��|@c�%��Rx:�T�C������>V.Z����=5��4?�9~�,ߥ�&�..;�yP/���r�R���C5��:��u �k\����!�����:F,�@4���cP��葌^�{�b̞��!�6<v���kB��K�ᨫ�aeN��b���M�'���s�oImJAR�R�5 d+��Y�b����[���#�� �U��2��H5X�ҕq!�Q��8�_"��շ@1v�f�%�U��aj������QMh=�R�����#j�c �Q����zl4h̗�=uˑR#:�O���9Y3�͠����ǿH���G�y}�{�97*n��~v/�!x�*5}p)�<J�7Tx�XYN���N���5�mΒ�OU}��1C�by�J"T��%Ik3-Ѷ��0��p�\Dp��_���-�)b�|�fS{��U{�O��@����͘�F�$9�8���Pn|�Ӝ1��r��k�>������4�O�ݙ�`m0���ʸn�ȟ?ز^u Q�$��Ъ��qZ� v�q�v�T��`�ۄ�,\Ӎ�����%�v�� �3(����Қ��wwV��捱�ӕ�����/���Z%�	��R�tKD��Úզ��s�j��"u0���機�1&�gW��W��^��O+"D��N���OD|�N��H��kƃPM�naH��ai x��r(Q
���"���9��8�_=�e�( ��Q�/]7�t΁ɜ�(��M���E�ut�?Ѹ��
8]� �b�y��в�XwBf�AXs�&l��i�~V���O]""��6��oh��*�~.��?�AMד�d�����p�>+��'�Z�AE���^o�.�;�I�:�ň���0�{z�^�%���|�c��[j*�c��/��@b��.���LuØ���{U��+tV�b(��22Twλa����w���7�&���2 O��U�G��}B���؋���?W�i�C���ޞ��-nM6T�6��{�*mM���/)'���p�.�oH-��FU	����_�4J�?�� 0휸��z��j�y6����{îX�D��`�����t�L%�e|=��N �[�@�Z�/��i�<�2�ύ���vyW����e9�� 	����ж�G��8qm?n��3k��o��$�ؾ��0^��l.v�ʂ,��p(���k�T��+%��^iu�Zh4�x�E�QL!����5�q��~l��=K�1�f�//�ma�T���*@����xK�=@���F�
�J�y�BjS��z݇eB�~^�	�F���(&�nfFqYj�U��ࠌ���i���?�*u�\�&w�cy���!��C��^�����x�:8��|�ݠV+Æ�����b��bc�7]+}��r��EZ�DJ�Gu�����5��׳|k��CW�HX��������:%�7,[?�)���0�$�V�;4����v�Mys��A�"�*YԢZb%R���t�s
�G�K�^q��F�,).�J�al��^�}�1�R�^Є:~Q����L� @�G�F�����M9E�o�"UI�>���eS3z�IAP���_��0�������3��(W��+r1�K��o�}��R�����\J&]8#4*G���>Ƴb~��81���-��G��v�ku�@�99F �Σ�%P=z7���K�I��ߝI:��T�֞R��e�A����/��AϨH��;����������SR:Tk�n)㄃j��O0�";��6yv�����Z=|�ߧy!��n��A�Z�9bwO��v��=Fa�ĥ�qk���"��Y��Ob��2�2�2G$19He�[���!Ij�n��5l�a ]P)q�#�rk�R���E�h�4xT�Æ��ǲw��13y+6���LTF0$�T�۸���k�Z#`y��F�u��c��A�ǩ�KeyR��W�+lA�j!���$|����4pDt�6J��q��ę)�k��l��Z�f����7wН����@������R���I�H�f�L'�܌gHש���Ӧ�k��%d �C0ǰ��ql��ٳ|�e;V5b��~I�gh��߰����rC�W�]I�7�O�d��_�X<
K�C�5��e����d����>k�]s�5a���kϢ=$�M2n$ԒȖ_C���v�5^���E��b�)h���v�A�|��>,����|(�`��̝.�yA�e�b�G$�*�B��h��
l�����8�3N�w��4?��ؠQp�#ҭ�鐨47�,Q�*':G�ǦLX�_Ϻ�5���5��e��L\k�����O`KR&lT�z�\	v�����8F���K�VE8V���9�J�8����d#��H��f����7�~S7�|anz��˥��V�x��Y�*Aк1��H	Y��̷��W�l�l�Tw��>g�'���_B���^p�O�I�����`Q �{{{/~h��b�}�]�aPcgT<.�G�l);g7���.��	�~�}|-��fT@�Cͣ���Tz-K;����l�[l��mU�cP*�-��Ei��\l�g�<����`�7�s5�?�]n2�����8�o^�e��¾�VC�NQ@A׺�B�;���#�l�+v��������t�!�@�>$	���,�C�<V������lbT��L(z�*x�ڻ�;$�zE�7��$����7�7�H�c\�H�5ҏ���(>�bK$�wԧj�yf�d���j>R����n"�)���2�eG"��N�d�VF=��K�X�-6�0��ߟ��� vH#Vk��!cDլ�6ػ��M��{���^���s-E��̪�i_�2�����Rvµ�@6c�#�u����W�� �,�O����:ב��#U]�U��t�W����j�'�vHB]�#z/�����7Ī�춦�ů����'��`�-F�oֵ�jH7D�R�":-..{"����������Oq,���87��E��R�p;�kqڏrN��n��s���q��g�����;2%�Z�x̧�bV�I��1�T��n-֝`-j�:�  Tq�޸�s@U[k�
ƍfn���â�F�L�f� "���\�}���5W*�t��>%0�K]� ��ŰG��G�f���4�qt@���I�������^Lt�a<�##a��b��5�]2p��ą9M#匄)��L-!wZ�|I��� �V�麂c2 ,^���:Td����^u�㼿m��6�@-�r������g<u��2U�r��Zkᐕ��5!~oiެ��PJ2�D'H�H�P���E�Pt��u���6���}�L*F]Y���gt��㸿 N~��%��������W���×�a��Gj*?��~�єk�4��@�uQ_��F����܅i𔭢�`�P��M�0��Y��*#��=�4�:+��f����YOU-AJr��Y�s�"
lձ_�X��H~Ǆ�&Ѡ��ȡ�>���s�A�� ����ǁ�r�F���l�IA(K�1�/��uP�w˅+	$��oC��/*IVv����ys�� *�:��y5��Ns��{E�p��'V3n�� i�*�9k�򠜸�^j^,
E �g�MC�0��L���s�P���9�ύ��=6p�u���"~�&KL���TZ�@�0%��/��y�#C�Z���£#� �^wZJ
4�7�lǿ�����:�!�q� ���u��Zhp��D�
T�iEE�a�j:��K��\�_�#O�<��5C?���Y��(0jܝI̕9�c���s��=!�AK���~�Gf�����4Y�x̂ll�M�U8'+��)Jb��&ưyz9<�w
�vײ9㛏^�7r�@y�����0`
�gNX�rj/g)�(�%-�Κ�S�Cb�E]�Tk �h&@!��T㚞��_YZ�Y�����H@�v�2_������������iu�ǌ����9�N��8���� !�mؿ4r�� XlxVHYEB    db34    23b0ͺ3Jx�D�����kB���"Tg~��1�޸oH󶜈|�8��:' ��\幔x.���i^�4�J!�׾���M�R� @�p�;�r�<�8�z{{���#wC!JJ@fU� �R��Y�~=e&�Ɠ�٩tI�G�`�\��*�.�^�>�؍�5H^�{���4Ǝ�ƠOT)G����+b��$���^��Qq�Z�jC����dTMK��|�-s ����w���8�if����V�΂���$G����-D��N�������S���;!�j�@2�*qD�L�O0����K$�{$�n��\�|	>]�KX�6���[�U��Ѭw���~�u
�y������~)��`!u����� �[� ��F�`��nҦ
?�&j���8V�Vd%F ��Zכ���(�`��$5�7�#��=aa�T�?���t���zW ��_�%����X?M��F��<��_~	�pk`���مP4ǃ3���@Vޫ@�����j)�
�[�/�odӗHiL�3���p���j\3cauT"W��͈��̱g�o�U��E�c>g:�ڒ}&`�����n������5��Xl�H���#����+�}d��8����F-ҙ�-�Z򟡓]`��衝���A���
�qkXIª}5Q��5K��"�چN��,�H���!�ON�p_�������/�GoK�]|薣P���l��ʹ���R�h�(��k�D��&�#XHw���}b3�F��5����İ7G�F_[��r8:Un^;B`�Խ��¼���͡�|L_��s;A�)�w��[7�d��N-�'E*��)�'�56�_��}���#ô6E��rm��^��3�]k��hĞ8��Q�bM�nq���z�z]��q_}ɾ$*�N�i�rAi�xq����O�sRt�z���� ͗`�b�a�(��������:�ßRks4ƀ�ʹR��en�aci�`nm���/��󎃌�k<=�����KH"�\Hy>t�;p����0�X�^Qg2�ޚ���?+���-��W��c\�!���XQ���P�����S m�u��`m�w���ڲw�_����ܼ�\����RW���K��k3�H��v$b-χ��!4Ң�0�}�,��qK��4�!��뻅Ň�wܽG׳Q�x�nKV�{�0fJ�*�~��~�e�ĸ��E�띱��g����������L���H���7,Ѳ�V�hDF�;���Ot���9,�@{`ܧ�"'n$����ѧ��,�޷�ME�3�$��A�!�)��2@b�V���CN���ݤ\��|S���Q��mh���G�T����u��k���n�b�wJ��5�;�*�����s���suy~�9�P���c�����KF���e��Ӡ�[ú�,���93G��V�6'^������ �`wK/��zc*���W`��	ȂM)x�G8AnTQD~pl����4� )M�V���,�k�q.U���������(�J%�� 椆l���k��$�⁨���*�4��]�}p�܀/�D������'�~k���UyD����������@�
e;��m4H3�7��ád��v���z_�@���C�1.(����f�*�)��k����O�j�@>��<"+�jMGX x>6ٌ�ٻ5����L����'����p�����m�dYn*4?R����#Ә�&��z%+�m��c���(���~� gr�:}pҼ�;^�iڸG�92�C��%B/N�|��|A������x�u��\��)�!�T-��y0f��p�_���v_��_(�85ˆ�zv5o3���m��h�&K$��Ūǁ�S?����>h��#���	�B�zS5��y�Cd�U�����#?����9��ZD�R7g�QëD_^>��{��X��U�;�����\��?�.�p>��<���t&��7�KX���9�ˊ��r���и2VDJO��:]X��A\�{�@ܒ �1�`�/#@�a"�_�ح'�N���U%ń�Ck2W{��:�����<���&/��0�aaX&�l�Ab ���Ov�B��V�=.y��c=�d][��%� ���	nI�|ǔ�Ѻ�9lx�I2��Қ�V���&���k�$?�pFL�c�&H�N��$�tH���Z�(j�0R�����gF[M5?�KI�P-$��h���[�PK�Uy� ��\)%�S��GX��L��ڗ�`�A��˥l����{��E���Gr�����t;%�F��y�V[U�NI��[�`�B�q!е�?�`O�����s|�[�_$����nL���� j�h9�8�'<���x�	b���<b�`���8u7�Y��=Eu� �@Ѣ�(�Z��PY���;��'�	\`���I �� "zGFՇO`��^�[o幈5�{V,N����V&K����'ើ3�ωO)����~�I����+ ��Yn��}y��L�K��a�qA��dU��{��;��7��tgY�/�.����@''�����X�[io�@�w�[b��f��h/X({A����@V�	���C�4�tΣ�C|�JJ��Qĸr�z8���Ј��] �H@���J	8�N��5�o#�nRx���	 nS�D�b�? }5t��w\y��8���ي$�хA�w��Ü=I�|r�O6�H�E����E�Ӳ���K���ǡ��٘j4ټ��ǰt{����n8?��A�3�E�0�a��a�n�.Ytc�T����0�-��Q$D�/T�fUQpASż�T�w,��X7��	�xu��w|�jmZ��U�P��n���~ҙ�i#oj�i�����m�1h�9��)5���'��t�,��������[��ۧ~�Z�P-[�f������Zab� �ߘm�Uy!uhA�m�3b֘�t�}�Ru��-���`%��:ٕ�?8�c���oL��NO�53&C�2��r�^ϞV����<�af���\!��U��zmVC�]�e?�}x��ފ�X(:Ym�� Z��7�}pJ+�.�iJ=;{��RW��>����=�(���i-��?�eDG6
�Z���{�f{�R��Q�n�*̘�9���A�t@3Y�h�8*����E@��^�	��?���Ė^<S*�i�l��H'�P������̞�H���
ٱm@Q��ܐ�xx��6����ln͹[��|T5��4;]���Æ�	%����%Mr����>�'cj��G�nf$�O|���e�i��s�����1�<�F�t
RX^p����i��b!1�'��@+9/l��G򄬓��Ժ�jx��?wx�w~���_�4��R�U3/�bm)U���R���5�������S�\��NEĠ�SO�'��z��+�S�a�.��*0V������۲�n7H������.�ӟ��T�#���mv��#k�	d42��YS61+��`8Y�&M=s&jC�_7���c�(	��gB�05Ȫ<)7ڟ�[	�9�����<��1����]��8.�lnS5yA�Z*x���B����%��/�b�e�J«=⯁�bLeɆ�T�'�R~E�\��c�\�{mx�ՃT���](�w�_z����Pꨴ���Z��
��5�TA��B&RM�1i��,�!��_�N��fK'e�

����Gk�68T�ԟ����ġl��V
<�1I�ο�fq�S��zgM����?���W��i�]N:u��l5&�5��w��!���S���fb5�{$<bu͔�˖?@O��S:A*�ɴ�wV�+���&F�O���y�y W����M��5�q���h6s���6��O��F����`��'W<�[ĩc�X��mmf�Ug�_�k��xM�ժT�}�\9A]�zr�7�d�W8b���;�/w�X���T�S��Z"F���F�~I�U�P¹]��qv�E\f���`�� 5!lG/0!�]��,���]@��� �
�̋�#������r�n� wo\ �:��{�����&���BPD���i#.�H�t]�A0k�vV3z[���d����mf<]/�cv&g��j�,a����w��H�)q|�Y��}Gټ����L�_�Kn��u-S�.cFKx`�ɩd&h8ޡ����l"g��T� �n�$ِ����Պ����I�Lڕ��.}�č�9�H8��>�7����i	��l*�Bvnu��� ��wxG�ƺ�7Q����V��Z)����].bI�����ThdNDb���=`�U��c�}+�Y���O����t��!\��L��9�Ò��y��x����wO0A�H��n?��a���jo��}�M�k�3]c�Tf�����oZ����MM�#�a��T+����&��\�g�F�`�v0i8a��^�	�ߧJN�x��Z�]��(�PS�X�tpI�ؽD�*�� WNI��1m��4���S�藴"��6�T٨S�/��x�I@�r����ֿ~���o��['@biC��L9�E��剄��c�P�E�j1�w���zsAΥm�[��Y&�:u�Zzy8]r�l� ��%���B'!|l�I��h�t��};b�V6h�EE�D���:S���8�2�zZ���팖G�N�/��@Ĭ9�0W��Α��i�MA;Yk��I����Po��}�$n���!1gw�D�"M~�]�ޮ�p����\[���E�V�
'���f����t�k�J2<���{�-�&�m��cQ&eZq���M�p��t�0�;�7�h��=9,���1X}�N�����.,�٧�u�}+is�ߑ7�9���d��	���t.q�)�c�Y�Ič����j����5@Բ��0̜���?|���J������ُ�#�!c�=ƢAE��O~h��v��c7�{�+@�6f�(�M���P�׵D\o'۫F��=o?!{'�dl,\������i��z[B�]���J2��Y�=��%�P2\�� �0%�4oU��}�t2�	b�����m��k�y�z6a]c��aaRj���������/3T�M���%��C^��\C28�2똪�ȷn��
��
��ɰ�7��s���UCү�8A�DL+)����P�T��a���ݽ6��$���v�JZ&��'>mT.�8����Q����{�����o~��2D�-ycs�O.s_�if��)�j��eNP�0E?	�/ ��v���0�(rF�9u�3�ƫ�4LEP7ծ�.�x��ڴC͜c'Jo��ֽa��w�������i�R��OY;j3��ړ,�:�j���I{)�߮y�ӣ?wR�{��O*�����r��2��q�˥�Lg�>l�?��\t�Z�]������E�7��N	h\Nyno���[m�6`�y��;p
���H����� o6����庩�m2wKSh�׉�
|�Z�kR�{u�u.�����c���>�ݩbEDH�4Y#��`O�h�3�
�I�P_�^\���	����
��MS�V��9������w�h��Us��W
^�2Dc��5y��~P`��\Ǥ�<�pK�y�9�1�`vA;TKY%�ǹ�3C�����'�������ոI]��x:�����U��}%�/���$z\�g[t�T���`+��BIi�*��	�6	������>��Ų���rzt{s�BU�}Nd*Moatm�An��1,�(K^\1bU��@� ��cq#$�܈���Έɺ$�JD�U�~[ݫ1�n�ĵ�<��R�ʢ�>q$2�|�u�j�!y�W���9�W�?����:�f����8n�j
E��X�k~r�S��GJ��'�v��%/��Ȋ	�'��������
�ƅ���M0�{B׃�d��M�|_ڞ[�ھ1�4�:�;fmv�d�v$�������y����W}a���Ho�v_��Cn4dmݜV��/�ۚJ�s��B{$�v����a�థG�e��^+��M�tw�#�\�'8�~���-df�%��`(��uʆ��2=ph�E���t�~��EǇ>�^ה�$����*���LK���믈� u�ީ+�׵!>�1i��t��u��(��͜��O;rsm�tc��R��������v�p(	����r�\iɟI2#�9Ď)g����h?�E�<qZ9`=/PSzjD��/E����Lx�T�	]����X.�)�i���kwg���4�F�ڊ����1T���,����#���uv?D��!G�SE�L�29��Z�hz��zC�򐔋%?N�!v�shY��c�;L�Y��ZA2໥W5׶C#}@m�}�[pڮ��Ro(�U�u�Cʌ3���ơi��w���0q���ks��f��;������k�ˏ�����a�js ���0CXJj�ٗ�w�f��+���PNMPR�Be	XGDX�ؒ(y]�M��XvǸ�F�*- ���u��9�fݴ854���nY��yB~d��U��[�j�k��E>���WӆI�)ߖ�^
PL2�= 븩�eM�|�։?��PYv4)�P\�H!7�F�b�8ˤ��&]x��~�0]�g��c1�D�	�G�G#72�
ډb�E�7�%����YT����P%{���A�OE�fu�ʭR���&qI�뎾=��o��� �}u��[<!D���c�Ii��z���9�6��%q���)�㹇&�}rzvc�q3�o ��㳐O
�[�g絩���6Y|�N�+dA����F�]�v�ȷ�<$�/P@P���b�[����WW���lui~ǫ'�h	g��w�'��=��M��"��rY�EU�"�#R��E
�C��c�y�3!;9�̼�u�P��5ęA����L�H��l��yw��x�Z&���«Q��
��v�)���;�b�Gt�2���'���@}|��^4�1����8���
;��B�i�2G�l3�ML�,7�%�b'y�3��"�I��B`�t��,��D���0��*³�Q�a�kb�AfLV�˦j3V6([�C�<�N� �9�O~I>��-ӳal���.6J�lz��1�>��*;��S�2Ω-���;>O�Ka,}F�k�+�u���c:��s�X.O�H�F��#�xл�#���m�����>V�M��~[`r��p��w0��MZ|�M��;3/�&������Fl������ψk9���U[�FAj�@{@����A~�=n��4L^�}{�M�K��a��C�G�b��U�=!��\S�Zٛg4�/|���D ����s��'�.D3�?�N��)�>������VK�.a��#��m�5=w��M6��9��7���,'�z��!�.LBW�i�l���S� �~�C��¬ ����pGGt���j���k�`�lل}�=B���d[=n}�,�_JD�0�K�ќ�J��� 8�u�L��0�<�4��e��nCy!��q�s����"��L��Z?�Z���^0O	@`�
kjKBW.oX��&�4QBC���0�.m(�:�7��<&
m�I4u�Tb_���A?���)N|��L���^�@Fh|���v�	N����6��c�ྲྀ{���m������hG��*�4�%KG���Hw�b�f��6��B8� G�����{�
#�}����f4|�Q���vRryFV�A��n�g+���q6�N�nڝ#�x���<G�CS��<KܦR>RE�L�heH�3�4.�i��ݨۻb��l���J.���B�M��<l�a)��x>q봿9�F�l�3A���VX��'9;���⟔{��Ɗ�H�z���
��-P�g>�����+&m���:�`H���,���k<
��X�,!�,�XhAB���4%���1򁽉�N����M�m��;6�^��Yz�1�\d���+��dO��ҿQ���ړ�_�U�q߸�M�TlV�vC�^��B!>�TJH	w�:���1��FJ��xT\ �V�W٤!<���-���2��h�D6 Q��Gw-�<�G�BlְCO�im�H��oe�ai,�Ŵ6O2ziB9nBn���a�h�?#����Ѝ�KX]5�KG`�&�����J��;=�n�x*^��q�Ѽ4	0�婇 �S���a�9ez1)�4O�j���;~������F�5�ūT��`���Z�+�
5��g>K�{˶�� ꁤv���m+�S��f�$ts�ȧ�Tݿ[[�b-�R�Me��e����Ҳ�vE��E����Vcr��m�!&���zBu<֡"T�2�<!G�S��s�u���L��5���j1e�j\�<�vU����s�Vu �����*�5��ڽ�
G�ZVt�8�ϵ]�1B~����]I~�E�"8� ,��7b�#d�^�s#�n}��\���ۂ�$�V��C,�يC�u�����^2j�]���*T��b@|+8E\�I?Cr��lX������-���J�\����
��=h�,�����C�}]��4�
�!������O���!ʻ����Ub5�?��W�E]��'�����}s��#<��U�Q�b��m�N4��p�����r`J%��ck�� ]K��+hs��գ[���[�Xw�>�;���b.��n&kVn��xV�+D%'"z��7�;�h������9e�Գ����Ё`Q��E7+�!�9��6q�{ܕ9�g��캴e>���Ԙ=r�C�?(�8AҳMi��ђY���ge֠w��Ǘ"�8�����|�|��8ۮ��~� ��-�_d+DN�pM G�B�I_c�_���) Q,im���s�{Qw��킾r���\j���$o�	��HP��o�>`�y9�v]��-���}[d�n�5F�(���r��n��I�a��Bb�����5龗�ʰ��l0j���uT��E��_t��_ #��z�j��<���V�5�^8#e�)����/�o�35�o��u	�l��{��k��o�]a �q�
F�N��N�r�J��{�H�<BF��Vьq�G�X{���Kc�o����0�Vm��v'�	ːB&�x%�l�l0�k�N��\�='���[ލ����1����j�