XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T,r�!��14�+-ʹ|/R�:��;;�zM�r��$�x�#m-n���˓ �?U�MX���D���t���?+R��&�uu����Rn�� i�ro}1�	���2�tQm�8`�b~o�B'�|��S��j2WO\`��P��ٔ%X�{���p^0���&�9��2�bgo�+F�clJ�ڗG����T����*7�����y"(�K�ؽ:
�㭃��W"_nf�X�U��	4�ȏ�=��j{I��Ѿ�d��6V�
Pw�(�}����nA�^�{�&�4����F��+ŇrB3JJ�D~���eP֔�X�nY�v�.�J���U�l��<56J؊��6�X.�@�C�:�����d#�A�ޛ���?���l���5�D�c[�K�s���Y�����Ϳ|1��X�͑o�C�Ʒ��}윰��R��7���ė>�Ui��V�:�){�g0n}�c�I�NPiP?�.T�#/8(��z�8D�����zlũ��U�,L�ޕl%��f�P6I»0v�0��I�(P�R���\-B�"�w�Osg��;D}@�P�菦nQ?�7�nlS$ �Q������%��l��/%t.aTь��+`�}WD �b�I�%���4�X�����dؗ�f���o$�9�ʢ�yf`��G�KtwtP�w���-�?��Y �)M}8s,;L��|4�����/����a�羽��#1P,LH��jWH��?$���@i����wn�tզ ƨ���\�Y}�'Cb�?�W<XlxVHYEB    5224    1740���������:?8�x=z��L�D��q!S��״�l|���WSZ�~��y��p��k����P\�&��$����rfq8�^^�]�� ~�W%�d(�C3��� i��6��Q�ȕޢ�hK1�����=�}VqY�2��[�?o(�����L�G;�3>�t�N�&\� 0�n����b��(�]�!~(���UFD�J��h@,�����!�\�����-�����w�U̕Ծ���^��"C��>)�>p~��{a(hu4�����d�0�,�R�#�OaP}PW�.�ZZ:��P(�ԹN�eZeѸh��<#��m�2'h�2T�_�
��m|�7X�U�d���(^��o�T��T�$X86��z�;��d*r$ƍ��!��::��="gM��Ut�ZyWHh$���Rp%k�s����Y_��-4t �y�Ő2��"!V�ٯ>e4Eē�%^В�+��M��v��բhn#5k7�8����[��Q���O��%��{�����D+�>�Ւa�p�ª̻�[��=\���5���`��
ϓ��������V/��H���
�h��́���|駾��� �3����ucT!����ݡ4��؃ #t����۲ّ�'�)k�6@�2)X��k��Y&��Z�Mh���^������g����k�s����6��:� G�%j��tM8�^�?{�_u��[Rh;���iG�:�6�C�q�3�5�I�"P�T}����`F�n��0&_��}z)tOH>{η�\��Liz}���`6v����S��~�5 \f2㌾:��?����X�l3�,(/D0"��U�����$B
z��=/�+ ��t��!�md�Ǌ�h�> ��ڒ}�~�秛^��g���,P��&y��B���jހ����]��W�Q��8��NOv�P�+\=�stc˒�3��Y#�%��=$� �5+_�� .I���gt��}��2��S�6 Ô�I�����Cu�l�²�և����~O4��hF�GN��b�a�s��]�~*��U��)hW�aO���t,C������O�r��%�s�;eJ�^C��BJB��%_?в��'l�V�M&߽A����J����S0�]7�_�zO�QuxH�Xѽ�g)��9�}wr��?Y�<��$�N��z`��������G'gz���q�]Od��R��8�����m{}Ϻbz����=�*�^[�	r�i�ɚ����*Ȣhت�u[�>�r�����:���(�m~ì8��%]1�s05�4TL(%9�0�+�<�͝�^����������b���A< &���NQ����\�
�Y���$Q���BM����p���1�Kw�\�i`���<��Җ|EёM�L>C�]hs6�F[$�_a��P@�S{��\�^(ɪ�2n��z �i�P��+ǾIẠ��4�D�Wڸ�T3��ְN�9������`3V��&uI
g�A�70�X�j�?6]��S�MQ����ĩ� O4M�+!�L��1]��xĲ�r�8wpyU ?]_]Q����8�VM�Q��?U���f?*�����2���2��Q_Z�L[��k����z�	�%|4V�n�LL���U~Kt7j��F7 E���F+��������a���1[{�ħ'��)U�l�T7��\�� Ȧ���0�bZKX��3Fd�Z�cW-�����s�nWg�ꇞ]����Xm}�ҹZ��9�^;s���-��,��M3�� ���7���%:�D)R뺬��ќI_'H_G�X���B�'@�B��4������{Tl�jbX;[c����ݏ�ǁ�Q@�sp*���G��ں��>�F�A�	�AD׻�;9�!S�7n0� Z�g�\��z���RS]C茶�i��,O��s�^k5�rAe�[�����d�%��X���F���1��R�T�6����-!4�?�U�e����|��˅R��g��y���t�E0��g]fǲ���۷�_��"a�x�s�`�#����ly��/gE7�Ȥ�D��=�c|�M���W��Fࡒ$#%n���ۭ����C���`���ܑ�8��05�nq�F��F��Jq�K$&z��C�9菏��c�J��N�h$S�X��2!���'ҩ,�8��fv_#����4�׸[�|F�S�Ι��r�@=l�ɵL���b��ɨ��lJ����*!s3jgֽ��Ue��kO՘������e�̢�������iΈ��7n���:�rd�Y
�]�F	����U�����!��7���n4h,4_�u������TH
ǩq�V�"����ɷ�9%�߮Ř�P�T�Q
��1�Z���2y�K%����ڒ�����^����1��֮�Ra.5��7��5�N�l��
�-]qa,l�G��ր���/WN��7>u��^��Ě��Z�T.Q��c�ȑu+�EqW]�y���i�8�Bg�(w�6�����h�K�;�B�G���>*W�+̂�
�9qn�����P��.��T��z-���vfz���8W��9&\"\��s6��c�90ָ+Zl-��O�͚(��K1՞c��'��9]�^��;�BY�:B|)/�y&��w�v���*p�
��}�гLY� ��SCm�й4D'G�Yy˶
�]�3�;8L(V�)c�׎@A����xtZ<�xc<��0�L��<�EH�H ܭ5T��hQEɰ�Ҥ��!B~A����X������.��9�VC����]��$�8�׎����-�'�]avׂ��dᛁ�ߛFhyh�p���crv�]�:$ԯ��(���%����C<K�����(�q��ެ9�?����M.�c�gQvEƈ�*�x��]`��`� N�4��^~2x�I)H�޿����ٰN����Pz1�����d��Ab)���1�4��T�r������$��r\.(��~\�"����6�T�
@�>�+W�U.���BFITIc>]\lf�A�U��S�ч�^�$�%��_E���o�J,W!(Ȝ�a�Y�ޡ��^�_�m��Y�2�@}$�(p��h5��G;�<��ѫ^Rh!s����M�by��/�P�$Q��h긟�]r�%��|��u�zj������N;cJtC���(�v'n�o<$�)����/zYv���� �q�S�|T�? N6�{ZEq�Z�"�t=�s}V��Mi�NƟ��u�^�6/���]�/��_���!�G�)�qS�Ț.��	�� ��tR��\��b��'�$[�}��gN[�؊�s�<7��� */.Ӥ25�d8~E��Hɿ.$�m)fD�0 �Z��գ�O� ލ���o�a�c��_���Ts�lTL��ţ@�P%�����g��ZU���ZW;L<2�����𶀐��L��Y����Q�#�U�k(�DF����g�W�x��>r��Iuil�3��Fqw�5��G�kuv0�塀xܑy��=�/���X����s-��"q������b��ۼ��:+�ӗ(K���u�HH/s�鱳�	ޗ)�}D�:5By/�C��U�x,A2���
�V㢏@psUX���
�ǉ:_�KZ��2�[E��ˬ�*��
�`���/=;aՊ9��Qa���j&��$o�"]�b4�ANT���De˺�}��)8��66Iy�T��>�`��t�C�gAկ:�M�ª�j%�H�y�d\EϹ�c�.�y�%�egA�tl��3*�\J����UQ�o�w	A���9�~x\�7�	vټ�Ox���-đ�3���j�����#����#y�"�%к���pp������KA�88u�	���'B����Su_�Bn%E&� mm��:<)�sx�l�ȥ���H̄��_��߇�I�H+iX%�a�&��4=ˊ�wI�L��4�E���ɂ��!�*~� ��7ߞ%!�v����t��� �LH+c{zI�:�ј#������Q����9�\��Dv�ˡN��t���Zi��@|����W=�c�j �J�@���z�tQ=�Q��"����>&&��4vu!�خ����Li�'gn��Өט�����:	TT���!�{4c�KD���&k�tm� {������\���>0}j�*������t `N
E.�i�M��� ��'e�G�VdX�s���6��ޒ�PO��@��E�f�2�+�y ���)��~�`�G���X�й;����wc��:RY�>d;�!���DԦ�?*�|�)��?}�W�)2�d��*#���{y�-����$�E7�������j�k5DR��1�&v<���m6����%u_��I�������:�`�$�u�q
��� �L��Ke�w�q�(�v���EW3vْ\��j	{٭���_�4V�Sy�^z:�++;+�)�mEN��i���|��6�X�7�vl� x�ގ�y;�h/M�!�)I�Xa��ߝ�_A����9���O��`�K>t�\&���ͫ3T�#�&�!�L�<q�^���\s���������ƌ��� ��/<).7�������e��R))͐fZ,������R/(��%^�l��x��h<M�ֵ�_9S�9�&B4�sT�@NH�xɞ_wI2�2�q�*���!o$w}�y2f�買�z�r�ζ���=;y�!���GP���8�j�5��' ��3n�ԡ�^%��@�����QsA��Eh�,��p|gCV���#����x(�����>�ϚR��X��5�n�e��1��1�Xy�灑�hL)��F)�pBN[����wv�M�Xg��m1(R��{���ڠH��&MIG@G��=5�07�d����L5ۍ�Z/s�BֳW���f�Ԓ�cJm�"�=��-��]/'�͐TW)/lV��G����f<��*���`�1����AS�|��EJs�Z�:��ﭔ1���ώ�A�uC���6,S���2ˉ��&����[t�IO�*�"\����Hgk��%W� P�������O�7����iJ�x����ױs���G� r�reR�F��U7lq�U�hM�0UJ�3��).;��Q�`G�	���$~B�V�4T$��h:�_��O�We]�:q)&�y�F�m=��K�������w��i���J� �
�G�������-�h����:����=���/)��S6FAdK{��ܕU�ÀA�}�CZQ%�h�ڛ�ߦ"����n����Y�U������Ro�ۭ2T֎<�3}x�����nou��q��hk��nC �2`�3��+F|+�'�]��@flU�}'�����T��E�<�G|�0�d8���eA��l$�zS
���w�kj)�@���%�b�����0�2"�AY�wv�z��D\��u�*'8<5N�d�\�ƹ�Z��>�GX�m�uyv�f��:�=>Ģ@��1��LIP+W�ѽ�5�);�gU��s�� ^�T�D��p�� ˲Nf�[�}��d2���us���BPq3�3��t���t�o� �w�Z~w1'�ѽ�aiU�H4�]�������7ϐ�/�Es��zx^:KY�wA���ԭ|�1�L��X�<8X��o�-�iqXW���=ɏp��=l��!+b��dg�Q�q��A*�V%g$Z6�L6U�o��JD����jbĂ�z��A��	�X�j�Y��C�%��:���WB��Y�]�j�u�3�����f4NB.��9�ɧ׿0\��4Y����\6�g�S���Z�Q�UL�j�%78*�哆���*���d�[�/lcQՠ���,�Q�,���(���p�-t�C�g�#��w4J0�M�Ԙd�T������P_�!���N~JuT4=OCuv�8!�Lx��:4i�_��'���&F���������sU�]��ȭ