XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=��B���M@�Io�KQ_�����N�������0�g�I����{1�,�=
,^vğ9Z���0[jpQ�,����B�~��8s�#ŷ������3y�a[����|�/��CRM�.�տ�#�-���4*��J="P1sCG�H��;m�kx@j���z4����=C��ѝ�y��KQ�%ym[ZBp�(��QƔ/�������Ǟ��ݯ�^28T��o���{>�:$n�)��z�/Q�}���r�Bye�ؿ�Tգ��h�U�έ�N.=Jͺ��r����_�u�����ۦ�Z	��ډ22���j����
��4����L����C���8��m�L��bv��^w���J�SYek�P��Ȏe�V��(�����%��0��Y��K~��ں�K��b�kd��ٽb#zxAv�߫*�*2���Z�N�$%�^tZ�,(e%�?��.JzJ�N��CmS��~k������::,�O;�����#��(��F&$8�*����l�1��|�Ik��x��x���$ob^�������	j��M[���3�Ki�w��OR��	��D!�Ivc��������XeCx\��RDٍ@^���,���QX�E��׼z��Id�9��?DF[aĴ�)IvZ\{���Ӹ�Yx�*0��DCOm}#~�0���m���=#D3Q�C�S�{t��j;-j�ӿ�͈o}ڧSVa���a̍�l+��/�����VO�f��ڀS?���m9�kW¤�S�P�3+�h�-t�XlxVHYEB    3e93    10b0~�������M�c2�l�գ�8��Vш tY� ��ڒ��F[F`�Ք<��rujܣ.�Q�R3U`D�e&�J�s^\�.ژ���r?B��Pgx�q�35q&!�}�=�}O�7]l�Q���|��j�$����tZ�=1�!�2Iތ�?���>�d��<�z@��������g5K5�0����)1��ag*d�v� G�i@E��|��UE��r�U�����3�
����Sq'qB�2[��9����2��7�3�>[�w1��!v����%��cۧL�FAQsI ��yb�8�Q@U��T���X^$�]7���O�x�*��ё�66��({���t�����I��X���N�a!�<�«������P:��G�Ս?l5�E�%�w]Pd��I��ކ�o�ꄚ5�L��k��h=e��~�>w�д����m�%�}w����Dޥq��}յ|B5�O�f~Mf�_�������?�kn�m�~5��L���
_��6o
t��
-L�pJ��%�`Np����b��,�Y���Pu�]�U��aej&NZ��	��M��{�Gt�l�g��J�MX���)��aN��OA3��}����7��� �o23&%��Jشsw@s�F7_Y�Q�=��n�����bT�ma	����g��r�?=k��7���f�dzvgX���
{�5M'�	��z�y[҆��(
�߇v���KU��5p27���NNJ,�kT~+���"��V���3��W�a4I���&I�b�4����5#]�mW�x���{��-"���o��ƍŶ+�*��n[����o�Fu, ��>��:N��+P�A\Z[�@4������YPw�/�-r�6�s�Z`b�<�1��.�"�ei�@Xe��:��Y~�*��O�(�o��Lo͜�~�����'B9j��}�Y�Q�~�M��t�b�D~��y�W�0N�D ����.�h�f�MW��M�e'I��|�i\<�+�!5+��?p���\�4*� �yU��0��s��i�b}^vl��Pn ㅯ�(n
���ٴ,R��$�쩇�x���
\p���9���B%�L�{D����#����w@�g�����;1�}����'~d�W*]}=Vhr�e�@Sl�/1B���\�z�b�:�}u#>Ԁ\=EI&	^Y3DL\ڮ�>1��}�ni9\r�O�����c�ݭ�����C"h")���ϼɓG�-p�;�¹��3�	g:{4�0�Ů��G�Gn��JT���
��Q���g�z����ү�8�3��0����t��iO#eų�.-�-֣��4	�X*$�RC<�J����@�0Nc:�/h��*'��}ʁ������R��J��|T2$�vpKW]�n�պ
����B�~W&h8��fT2�P�Y��;�����|?�X�m\�)��d���U��.�)FƋ�$;��~.��JPa��rƇ�k����J�~��[!_�r	/�^�>���%��X��\S��j�?ݳ�'���)��
�V���B���aJ,P\CF;����;�{��P��0!�ya�6D5�]�4j�Tݪ��el�����_YK򫮍��`K̿}d��y	�����I���̿��E+a����^�J���R��G���s@�T��;�?�jv�.��[}G���5R<�SԬ���0�n��bZ�����L*� ]_�[��n�PDK����[�&�T�j�(�P�Y���~^Dy{K*��Qt�q����x��N��r��G.4������p���wt($�턢����2�+J�� �ҳ�$j����x�l�&Nz�*=�\�à\�x�9.���O�I&]UЕ�>�S�4���I���M��L'��?�ڡ�p���8t�a� ����]���]�jk�P�"�R} �jN�,Ø�'�.�0R�*���I��rg!�:���/>�����.�T�C>�4n�+��X��B?	�a*�d	7<�<��s�t������d�2CJS�B%oyzHJ�3M�X�qwQ8��|���lGdd
9��T�0����9u�p��$�#>)9�#)$�u.W�R7�Y���e ���� ���mb��D J󀪕�;;dE�cҐH��X��x�1������>�1�_ӗ�]�,M��r^{���ʂӇy��N�ЮY1^Pܛʬ8��$嬈���(��)�t��VD��!(A.����E{7�蹡k.氒d� ΕxK���K?HŘ�H\��E��uԕ�y%�=l���&����ͅ�n]���E�WG�%��3�S^|�	����c��JN+-��K8��K�����0�����niO�$^'��UD���E��k.�Ls,Ї��0R?O�/As������Q� O�d��0aDB�����@29G��E>��ɰ��i��jiG��:x�*�J?�M�U��h9�dCjJw�(� ]���݄�>gDz�;�Lg�v��P�4�=��w��C�e0<�M����a�}% ��'L�����:���R,Q����B�U����F��ôm?T�±�q���d@�Yئ�����,���J]�xjt�ؙ�ND	�[�p���c�a�����υ.)[:p�2����۽͋�/]�&���f-�ƁC<a�i�F����υ^���r�2������AO������R�&�i��P����n�"���C/LT"@gC`]V�5y�x��1T���0Oe���ԗO�I%H�8��d��q�v�z���C8So�7���LWv(�3g�ALP��յ���B�˗�fǝ�Ĕ�f>g^���Ͳ��_&@wM�hh������KdZ��tU�E?46�PqV��q}ˢ�����5��Q���襭�l��������nt�`��i�*�~!�"��
�k���\�2�5��RW�9�N5*�g�H6H�KG���sD(���Bߐ�����)���Ji
Н5*���
�ˇ;Qr����dr܍J��Xb�=�ï����xd�֧�s�o��L��˴Z%��oP���ď�hҬsZ�D�f�
�|E��K>t��U����hjbF��4nkA�H!ܧ��
Ș�Uf�t{�P\P1{H&Y����[�q ��L�3%�4���Z������5���{����{ ����0��������(�zk0��k�j`wʁ���:�s����/���_Ǚ�@#u�
Y�	 ��T|
�T���D�gb�b���#y{���km?����m@�|�@ ���B.���vD�uG��oPQ�����$E��L����7��m�l
o+��^55�s��%�L$v�E��%KP4��,
�8�$D�r���/r�Vń��b��ʷ� !w6ľ+n%�(�w�݆o5|r�ǣ[z[f��s���ҋ)����0��(\�`������ʯ��I��=.��r)�YDv�'2�/I�!�S�-�'�L�P��ڄ� {�x�>cK��1ZGY�������H�k/��%�E^(\��	�	uh�Pv��d���h�Ʒ;MŰ��Lv��l��9����i�$�+�����ib5�DF%����\�#�h���S�.�=c�]jT5�
�\I��������0��$��ѧ|Xw���>������?YnєmV4S�CA~ﳂ�`x�����}\R�����B�j^-L*bR��ON�R��5"���8��E��{�S�G�U�)P�w;N���0�R��4��WW��U��Z��*T�8������y��s����j{q�rv�tIm�E��4K�F�uڛ���}u���I��C ��6L���츍������X��a�
�oF���Q�Sڽf�./�)����&�%5�&ٿ�'�c"�*[��l���N<G�>�u�scA�䥪�R�rtR�v��X�z
	��:�PczdFO��E�;����_ ?���3�H~��	���Of-��m�PM�PG��	xL�Rl)���pqL��|h٤i����Ǆ>T��wh�-���xr�֞�F)�Tn��h��Y�7�55ϖ�i����bu[(�����g ��H�[2�ڨΠ\V� ��acӷ���=�dM�^��m�>`�B^�t4@��%�O�ч���	fc}��ׁ�������q}H�drG����r�f�a�p8nt���eV1����<P��j�8wz�&�����kL+�L