XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���&1<l�6��^m�ݚ{���z�Ԫ[�D+��յ	�%�H�~fY�_��.�S��2t8|�&�_����½�5�/���-��-M�P�H;T9��Q �o�){�)!�H_u|V��m$���6�������I���r&�J1@(�og@z���iNЗ����B�N�F�V�%�^�ر�_�q�d�lYN:8�T�5*�wE���q���������Ug�:!����ӛ�$�؂筜�����Hy/�V�QE�({G��w_�;ؼT���D���W�-�9��Hd�d ?�2���L8�C���~�<��B����:B�~RZ�W����(�.D?�"	���O�T��Vͼs�����Ȑ�?9Y��0JJ��p�������*��?��e�Mn��g�S���m�)�]�-�V���vJ���DaH>l-�㸠��Hy�L�9�4���Ip�5�f�n#%���e��o��İ���o	+� Q���Q�A���m3��8}���(V��`���OD�9o��su�u� Lf�p-3
�ӣ��x�h=C��R+��8|�\{G
^�X�����t恝�ج��{�eB�H�3�������~���/lK$/�*Q�Ko����E���,�y�C��[�xE��G�p͞�>����7y{��Wk���){�4M�::q��G7V�0�����I�sP01����+1�5r�.��-���d�f��G|�̫!]<�{�I�HN o��^�x�9���"�46:��h6�4�P���XlxVHYEB    39de    1170c�bD )}��ao���̂a-�ꎚG�EGL�c3�"�C�H%AG�,�{0�J>X�B�t�s�\�m(�!1�O�_3WC�C{e��"-> i��ԪPOk�/����T40��C��쇍�$���[�ɻJ�>=i�hg���&�q���x�����i�B�0@#��W�D��:�� gBE"��k���Y�A�C�nJ,0h�za.�Oh����A�9��˥��Gqu��{��˨��#�c�n��Gs`�^0�$5����7*'1x�%Q�vyW� 0�؁[6cr�	%^�3���t�L������!~��0i�
�;�5�,qW�Œ�D�SȮ<F|�%���7��Nڐ�4����"jŁ8�X�/�y怖"��ld6k߇/��rG��5���'7S��|��n�L�����}�
�V�r�l�#������\�6Ɨd��u9�S\�r�H�}��X�E68��6�2wۮ(�w�=5@D�����1I
��y��[�������
�p�gtcv
�K<}%(���1߾�s���u��KԳ�:�s�+�m��a��ab��á���t����Z����T5���ܱr3Sի9���z
���q^Ns��\,h�W��*��%�(`�2���<ȾR�7q��-����pơ|p����O8�����e�x����9��}�i�^�����u;��s&e�ߩjX��{ �k1l�6�����K�d��"/'�pI�A��7�y'o������?ԩ�x=��/-�*�l�L֫��G2v���ML�r�L\�97�S���]֑��q:��z��@r�i�?�dsȞ�B�H����#�l�|]��P�ީ�(�peGjy?��#	�[0j��#I/
s�:�K���rN�WUi����QCz�\ћ�k:��υY�D���\2�i�r�L%5<<���=$|�L.^Ɓ=ʘi�hc�]a�����ɏ6��sT�e�^f��Riꜵ�xZ�����������yWh}����Y�sp>V����{�cy�� D�2Nf��3 F��$}�%TnU�Ⱦ!�h#��2�5.��|�Z�&O�Yr����>�kc��m$&���U/��Ћ2���77��VH,7���4$)���.Q��M�3e>,��s��T��������iu��&9_w���ݯ��`c��,�ɡ@�x:qJ�磳��#І��I�v����U���!���j�Z����]�N,��i]I�#�\���s�3uV(�-rʏ��m��K�b�%���V1�&
���t�^�v��j�^�@_Ǚ���+����%'���O]JQ�!�OI֊J��*'C�o0Lx�%�H��?a ��U-���0Nߔ �A������o�w���$���if�#�9fTn�ģnĈ�H����&�x
~��u�d^��g2�/mf�$UnB̙�����0�����rы���3�p���я��]��,y%�{�:�kģʿIO��F��m�u���@w�9��=�\��!�q7�����F��\q"��������@K6Ƞ��9��,A6#N*KǢM��k[2�tTQD{KK�������ޗ�֎Ǵ�DY*�g�I9�? ȉ
�
��$3�]�.eAǋ��n7���,��<$�!�.�y��>�AiH��̓�Â�x�BdT+�3+S��.�|%UR7��A���.a��{�&2�W����`���~V<��:�,h��-}����M?��l���'#{`�E�f}�G��{�4���߇X��(��a�+�ҭ���˝�����ܡs|\�Osυ3����5�r~�P��m-���(��s�i���^{�X��A&�]я�j�y���d��%��J;��Q	�,'�i2�����Gi�F��M�������� ���:���;������54�,Z՟�Ī�t���b�[�ȴp��2�o���x�s2�����ZB5R�ͿEpW)��K���,�18�[��N�ɫQtl�!��i���O�.0ک�B���H^�S��i��U'��Dg)X�8H���%��ٗ!1����yԨI	��Q������ZC>�e�r��Ձ��h��8���~�(KI�(��f�q��'�Mo58������g��R�����F.١� p댏��>���>�`Q�"��Y�ߒ,[u�Z���K*v�
C�ToDf6$��EP�W�'��� !H�#�M<Z��zB�n�vX0t��.|WAI�g0сbYh�G|"VgRP���(Wb}AЈ�*4�d�_ƹn�@5���<�ȇd�Q�썑�����P�E4,���6_�;� )k�b���r�����oRwwXY�/E`*�K�n�&%a�R]��}�<�����D��JsȎ����2MSVyo�ȅ��f�N��Ȭw�rm����R��6Y�5n���B�(����:����8��K}ī{��ɽ�V��ڄ��������3N�-�'Ekb8a�2i��ѣ�Umm������j�Ot�1�C�c��a	jPc�e��T+UwNq>�ղ�!fF9�L�'� �
)��0����U{V�؎�&!&���������pP��kP�9=]��-�cHCH� ε���Y��K!��^A|��tI�Y3�eۗ�S��
��[eE�ZF�7�YL;���\s&m;kNHNv�PΝ^��'�<�WB�N�?� '�h
Oo����#m�L�{%<4��/Ȩ|�ѬbE��H��c��'��������w������;s��	�{�p�4�Q$�o��������'Q�ϖ���7kƛcxI�����t�#��n:�˔<%L�N?ŉ.�?�?���Ιv,�"%!��N��s=�DT��s��A#�~�=Ӽ�,�>s�ɬ沮���Z��%I寡��7ը(�	`�\��[�Iܮu)��B�o�(��[Z�O�{G��a��m�"xv���"��:���׊2�����XM���W� a��t�]!A��ڞN��S%�-}�5�kl�8j�`i�d�̥"��{C-����������sє|1���(��O�3�xQV/�]�f�v���~�s�MyӰ��wE���т>k�
��,�����/<�+�=$qɃaE�$�i��W)��O�;�9��tw墈���,�I٧��6� �eX��^��H��7�����ɺ/����f頙H)�
��:8��`�.U=�r��6}d.�ReҜ���)�S
i��}�y�K����gې��Shy�U�x���1Ԯn��i���|��� ����ݶ��ӿݺ-�ǽRo�!�mz��ﯞ]�b�<�h��w �'�u4��B�!z��"mQy�b�:�VN�}�Mj�?.0�?6�� �2WV��z�)��ٞ�l(s���zY�~l��6��uj�RߝeVi\i�K�>�w���� �i��[ͼׯ���
���4��Kx�|~�3��R�Ӄ8i��!p�z�^�w��,�Ә@��T�ֵ��)�z��g09|v����iE"��zHX��	�� ��$a���nҨ��}e2̕�To|�d/xɞ-6����+Tx_�sմ!%/G�F/y΍`�
�1KN�I'�QvW���[�,�)�q���@20;�L�H�%%;U�� ��S�m�Of���选�p�R�X�9�@�=��������,R�;⩏!�m���s}7)!o������Ǟ����fT��^��m1@TS\�4��VD���[es� ��\7�T���r�jV�L��=nc�Ұ��c=w�(�����d,�d,���[%��Y7��H�M���r��@�B�*���h�.�8M���eHáot�$m�mp��#�d�gWߢU`���j��/l
Z&����V�����G9�� ��lz��ԑg
iQ�*_a���泠ڴ^`T��Sc�V 3n�܂�А�2�7��[^����(�zl�`�9�OD8 ߎ9��˶���1�k�MmTO�@��<�,T���lG@G�v��FK�!#E�[uB沈΢�qX��a*�����)Aj��Ҷ��W`��/�����@���sc���'+�Q������ /X4���ƺ�K {��Jj��D��
�Z,4[�1���3�� ��2��y���2r��yߒ��U���;��,WeS#�ۤ7���g�vI�S3�i�e!���������axJE)�]X�Dr�;Ө}��f����4����0 |Z���SP�����/�毐|�����N�j��̖tg�KT_h�#_7�$`hڂ�K�����&w���wu>�T�
��Q�`{����M�CL7]"�������nς3�$�z�WP��9*H���9zP%*��RD��j-�{K��)�$�${�p9��0~�"�Fq?BOJ��r���� ���� �%#9��� �\���m