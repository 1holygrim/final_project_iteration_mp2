XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u ���靮\q���W�Ee7���M�L�R�%������{8<W�N�\�I= ��Oj�;�͓>Tk����� �U��!�ѩy�̆��'Tr��_�����.�f ��!/i�=���gEO3����*���oZ7�I��˵RjaF���V4>���ou�H���`|��M��1`ې(��6�!��g{C�r�|N���T���㾀hHzs�\���a���.׫lѹ��|����X��Z|2�E7W�U^��#�M��pm
`�^�_���T��7qV<2�Zm)�ٝ|=���r��b����hv;�ӻ���ܨ��3%0rܫ���LA�D���o��"�j�?=,Ib*n���xV*�o��%p�%\��9���K$}�S4N��7}x!=ۡ�`��4`���r�����K=ߠl)$��$�9+~�O;�9�՚ͮ�J0*�npB��'��l]n��[�c�f9֍�'��S�F��	�-m���eV�4!�M���x,R86,��(���L-K�HxAc�Im�^���j~Lb�~�.ە!+���<��3��Đ!�$�{^l����5�_�n�l�`�$[F�l� چ9LMRq/EЧˀ2���nG�t���N�����=*?�r�%��&��b Γ*���w�R�t�P��G_��G�}e�kO��`9��!hu������G���TfS\��%��pUb�s Ɵ>���|��߽c���C�l�@�Q�ug��WSn~3Ͷ���AKh5<��f��XlxVHYEB    1853     810ʇ�c�[I��hz%��Z:��Â[�R�,�!��^CaO������g����B� G��J�}�K�S��-6�I��P��J�VK&R7_6�.Y�h�3�`a�:�2���Ӄe}��G��'�4�I�?�*(��4%:�����]G?p%��D5���{=s�4���`����p�; ���3��z��
��r#���D��!�}6����4mZd���e���;��e^Z-����s��F�6���)AS�ΊfZ,��(r&{c'Y�\
�WG}�TFcG ܻ��S�|J�����J��"\�cO�V>@�\;�ЍA\��5I�^�B����y��%���������^ctfD��w����Xj�jxAi�
Z�����M�����bJ���9!z�R�l�:D�<��RU��]�%W�1�/S��_tG&g��h�Td���]�c�~�s��O��N�.a��pV
��w���$�����Â.�WeX ��H���>=h}��,b9�8�|}�p\���[�L���Zg����7��s`@��1쫌¢
�5�FM	����"Q-�}�实@M3�T��X�.��Fu&��(u��$����)J���T>��Ko�g���,����v�P?��怅�4�,w��o^	� ��u i>JgB!H��=wbؒ:�\�=�����gz���6�ttGM������|�2L������$JD� iDz��j�iޜdjzl��E�d:��T|S��}d�Og��f�f�?e��B�ԃ?8����m��ޢ�� ,1��Cԓ߉4�M����X�ђ�iqi�L#�ڏ@O���/ڒ��i�G�4򏤴�:=z�O^���մ�eZ�ʥ��+�b[���G_��/\q��u������g"{�
6O&�`E[`s���ҶV���'���y��7�/�O�� P
��{(F�Έ��'DT��Z|��U�q�4)F�� |s��/ע;� �����~Q}e5�Rͷ.=�'��+t��j�H�T���,���.�T�>�n�1���W��-��������Χ���*� ׷B:3�R�Ğ�IT���[���Z�2D1������_�1<Qiz�|�R�� F�>��T��v<w���q�"Y���NZ�Ę)�����hF'���>0(��f�V���Aӭ��+Y�
'I2���	��nw��s1F��R������Ubhn���U�1?�c���S�-�,�(�IP�Z~;ߠ�d>蚸����x��T����+�4�$&Cێi�ᓦ�s�9�b/,^*�0!���\��"�&����˓��΀vl l���9&;���ı?�R8��W,/�����38�[��ɟ&��+2b��ɢ�T��1n��E�m���4+�Zk��	]��}p�D�K��վ�gj4��@��Q��z� �4������2ReD��ꂋv�4��P_kas������C��^@S���L?�4p���2��u��'5b�͜�/����v�M����O�}l�����B�%+����G���0��2�H�)���ﲣzJ���Ԫ�a�z��g�*���qf��ДV&3���;qa�����H�����"��z(��U J�w�v�uRP6���>�g����YQ�(B�r�;2�e��ˮ�1X/V���+��z%jJݵV�l�=S�o��z�X kw���˸D��ϩ^y�px�;�2��V$X�fJ�v�NJ�öp�2��<,$y趮 ���K}���_�D��.� Ft!�8����.ī=���i�){BށÅs�]e�䮗_����Y� �ZǛ_�%���eLw��"����f¯΀���'E��]������-�,!�D�0~g_a��h*"��S!`�gv6	�y��k-;W;��g��?�B��=�jԇ��T�5��m�ڔ���M�*�|�=�g1�8�"����n8�u?�m#��� AZj�@���^��DH��V)1qq̼܇d�7�SqW���Wf���ss�����V"��fh���"�b�QC��9m�ĥ��=uP�@�񱍯x