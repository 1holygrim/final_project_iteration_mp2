XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_Mֹj���~ٌ�����x~��˔�᧾n5�5�g�X��i��8� H���R�?;��5����Zsް�N�t/6xdx2�����+��}��4r�R@L}r���x_��#ۛ|~nU����F�}�>�?���V׽�K����¬��h��4�YZ�-M?NC��'��}j�P�w��X2��*ڀ^T��d��D�Y��c��썜+�r~���@�!�G�(���Xy�O��!B^֡�i�l��֏���`@���]:d�C��Ɋ����*2m���b�vv&q�j�\&��m/�6�܁��Z���c�f�'[�$�'�ӂ�
�鵵�
=+i�x��l�q���ȽWx�m7�;�׻��2�'�-D6i�M,f�/�1�n�O
�;��#�k�B���;e�Ô����� 8w��4�8��Ѐ��N�d����]v]ٮ�n(�t�a��> xNE�U\�w��B`?S��e��)`H��F�|xh�f�.-J�9��M��+�Rr��c>���S��-	:iI�����[+nW�P��_#��/�M����bNۥ��^0��9�L���s�֠�$��G��&ͼfG��2s�QyA*�	��DV�l��o�J��]��H��x��|#���r��KC3�kn���x���KQSw�=҉G(>]EF��p�剭Ny����#)`@̇f��q�����{���9��������L�v�#��E�Ih]iBcL ���|L��k)m�f:���Z��eI
ڶ�4XlxVHYEB    6653    10c0{�'�}�ږ����aZo	E*N?��폿)��1ˊ�a?�v���]�j�e`�ѝ����_{��u����y����.g%�L�b�k7�P[/�l�J���Lj�͑�����|!�2Q�ŴL�iT�g(ƲY�f"��%`a{�[w˶X���)xj�2x�5�'n	��a6�=�_�EʻR��DB�m��)xH@�*+X��Y3���P=�PY��Z� �	��^/�-1~�c�>{��Z�;���ue�//g��}��Q^���bs$͔ڛ�<�ҝ�p��'����x�
�	N��X7RC�ϛZoV�������g�	�4�G����%_��w�5!�dAǲԺgiS��l�/� �=Q��C]5��+��r2!$T|*�ҍOTƦ����껻L�^�)�
�q�@���-�}��`��8P�Q�%�?'o�qI����1HE� T$���Z�i}V�b8��g�������s�{�J��t�,��\�k�2���Q�0��ySu	S%�S���l����0ҥ��p��Sd̙���g�d�6��� $>c��V�۞p� n�1NHT�}o+��y�4D�Zvo�l?
m2�[��}T��Ǒ
x-.J,���c�tzF��7o�W��G�Wt[^��n���Iɻ�tS6�;���ggAD��u�瘦�`z����!p�8��g������8�B�Q����B|J��{Z�o� ��s=Dt���O-�b�����=��1����B�yd�k�E�/�V��m� �~���7���U��B���!��x�Ⱦ IFc+\���%a��8/�m��p�D�e�猃d.�d���Łm�-0�i��al�"k�����9$���-�5� D���=����sʍ��P��.㒲)r:�@/HX^��o�o�3;���Oq��N��J?�1԰�����2��I������v`��az�r`9'�=��W�V�o��ݤ��%�Vɉ;�L���pk^N���>l��WTo�u�U{��$��Mt�e�.��u��|�A���:m��VA�{�S�'4E#��-���kx-��n��D���-����]C3���x���;,,��sE�p�����_���!%�|r[�݅���YY�~ţ�������+Žd,K��NLg��tr�9�a��H�����6�X�� �ʖ��
A�bԬ�ʏdď|j؟�"v�)c]^�&�9$�~g'@d�5"�u"��Xd���|� }��Ԩ����E��-6���!��L�@�=H�,�2l
Σ�cQ:2z�w�@� �%ݬ��3��V�K���&�m�����X"JW��u69﹫8t�7-2A]���N�4c>�ts����}"F={e%��/��� 
0R��הB84��*����N��By��J3�s�����Ϳ���-#|d�LN��n�1]<�N���k���cܙae�('.�#��� ��m싘B��z~0��*>xCP*�&�V��"E��Z��� <�xEF�'�3r�d�,%��]P�j&��`���=�3fD��=�k%蒙��2���z�k�qٽ� \Xiڲz���J�H��-�L)���2��4i�Or��͍[�����z��9)5�>:�{�2g����Y���y|�N~j�n8������/���	�u��	hy�ZmeQQ�^G3bָ�&�H���nJ{���L\;���;�Ӛ���Rk��l�S͇%$�{��E���|}���e�>tZ�� En�r)X����e�U��2���)�E���ԧ���D��;��I�|��Y��l��>~�.�j�t�㨴���e?�*�&󓛘=��샻�z��{�oZ�f�|�Y����f��� ���n�6/n3��!K��/q�{[�=Qv�-x>��7��"�'�^��H����
�U�Զl�h�lē���t�j�u��B=t���
���>�񕴬�Rx��'�Ǒ�,~��~��O��3O��J�i�Bs�Y$@G7��ی���}�������{q��'�i��"����YM�P��<�m8��9���Qtһ�����V%�.��<H��je��f�j�a�#�;7�@�b��eGR��b	�]����$K<"��Ê&��σ){��<@�����ٶ���N�K��<C�e��6�᳞BU�Zt[:>�6�d��x��q�AiÈ�S�g3�K~W�>S������/���Mrܰ�a�t�����;E�s��x���Md���J*m.~p����-D(W_��a�+���k����OB-HL����8|��&sV�ʃ��u��D'�y�A��x�U��]��{�K
$�׆|�[��c���C^�ЏMѫ�j��T�'���K�:&�I ��g=��TC��/<��U��ܙ{8X"@W[�����h�T[��r�<�0�g�m�k�#5�=?�m��z�ӢoM�kVq��\Ba +)sZ����Av�KU��~-���m���;�at�x�bلhֻ4h ?;iK��%h*����T�{E;�H��;�q�����Qv׀ �n5�u�;�P��$H���BF����R��zj�_+q�u�x��\K���Ivr(}"��H�T�X�p��S���D�|��eq��#����~>���p�m�!0x�d�4v�-�`�x���>�.�ώOհ]+���Uv��'rUD+R�F�3��,6d�.�~�F6ȇIyH��񨋌�C{}��Ny������0i�ڹ�X���/���Ł�:I�l((Sű&Fl�lb]��?b��	��W\�U�"�[#�Pfۡn����E����V�=�h��<w���g��B3Öx�R��ΖMF���3fCh����`�
WzXfX��.�; �U#2�V�_�S��Nvu�Xg�[DJ�1-��Sv�X<��{1��B/|��\��]��0���/kw�U
Q�����y����j�ue���7~�G]���H��' �"����?�c�}�:CB���k���1��N�L��n�q��^��.�!�[Бi�Ր�� ��Jر���i��@�$��sW�|�#wJ;��fJsGB&��oD`17���n~��d��(�v�]Oͻz�s\�'to~gi���
냢����,\��x�H<���Cb�d��O'pk��J^
9tI6r���=(��x���o�f�m��{�}QeQ��+���9�m�*���Cԉ7v�:#��W�O�ށ�¥�k�l*����AZ6�
�� }��*T�܁ϭzt�^�8^��g������U94;�!���2(hx�ק|#��=y�{B�G�H8�C8a` ����&���~-�&p��keg���'i���λ�|DR��)�j^lэv0�?��P�ȑ'A�U�oy�hj,��=\̇��˻��7)�|A�`�`��8j\l�%#��������ݟ�3� �M�O8Cq.~��w<-Sn�!J�H2�̉<ϥ^��A�5��K��37�UqCw�m��O��7(��he�
@HXI⯺��)�)��c�_�Uwb�S  ���jp'П91/��!cj��TR��Z�t�A��b�J�%&�� @7������)|���3AO5�_E _���)��#5}Ua��OYf�ʑ:��E-�냇:OM��feQ��iK��E�=�=���G�v��}���ma�����y��숅���Y2�K�7���=���+���^�4��e������3��8ɸ�.�MYϽ=朹3�T.s��L��5JY9яD�ќrAk�uy���/BC���ue>se�sT(��P9O����{Y0�	��f�"���{J�T���{(jV�Ѧ`C=p�:e��8�uɜP�P�n�3�M�y��0����`逰��3>l��\rM��L��7��P-O�'��62�V�9�!��e�$RZҺ��@/s~ט��?9��s{|*p`�i��)�]��	�ǖ��Z��R�O��!Qg����W�JʦA�O��^N�J�^���fE�f�k�=����,��g؃	>6��*%$'w���kQ��_��:���z�.�T��GY�>uVs�O��'v	���V��o+HȜ��������NJ|������&'���#�zO��Gz�̼S#:1�t�?2d� �t@�hA8�v�W��R�Fd+��Dq���������n���0�D!ҳ�/�����Ng�pw��R��Շ�7�+�