XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E��b�a����� *[�Xo��]�Kӊg�,̝`�v�L�o�e�PJuA m��.)Ab�SQ�_�,8�}��L�5ٗ)�u
�ժ�#��ϱ_dD,n�ȁ�Y���k4넴a%�%�_�y4=q�N�3�yK!�о�x^�9�ӕ��$%���	(n��lz��N60+����@	�t�mF�l]��8�w���$�ӑ�"~8D������^�bE�]�s�G��e\��It%l�L�ES�a���l]z�L�mG(��F�k��CՐ;��؄|t���8�ݟ�WX�o��$+Z��6@����KM����?sSa��@(K��ڃ���Ȩ|� �g�7[���a�C��(�mM Qa��i��+K
�t��D[4\��3ޟ��@E�)���ǰ�3� ^����ֱ�o�(c����_����ܽ��ϯ;J��O�3�L� O�{�z\�U"*�15��?��;����$�"���\SSN�LS�샐��@hxľ6N�-��ZY�ej�)�)�C��KFX��*XF�閸�B��V�>+�߼�@
}D`�T0M��0���`�.�q=�Q����y˘��-�_������� ����Wd2�C�ʵ�MIe�`G������r�N�����/�N��Q�9'>��ϴ��Z�z#1�~�����Z�B������-��B�4�jI�<'J�&3O�Hw#�L�\�/�(k��v�#�/��/���M�p�L�j�[�ċ9�.6A�O=��?%��uL�m��]Q�g�Bv@�XlxVHYEB    da59    2e3059Ũ���3�H��'fʘ����*���mr����S(���2�t!]lS��;����Lr�j��4�y���>��n~����A�͓)��^[ZG�˻G@�RZS��[�!�_a��4��A�q����\|��P��3�m��,��:xz3���#�@E������Q�����<� �b�D��.joX�Ω�<��C�:�C��]��5sϯJr.ĽE(�W4&�P��������l�3�����93�>'=c�d���v��B���	a�h2��۪f�"���?h���f��,�_��Ji@y6���M�D�@5K�dSJ�}��.�����
''�� 2�!��Ƅs'
����"��܅.�6�jO�w�&�t���6�(GP���E�f��K5.�9^�(�N%qWRa�h\��0>yZ�#���
����Y��ʋI,\?J돕���p���P�^g���C�D�� ؍��>��/����+uS���+�M�B�WT�u��ۏ-�Ʌ��Im��s�������<˥�A��9ΰ۲�E�m�fq�5�-3]��>l �b�X� Ӊ:_��T�a��6_R!�
<w\H�Z��Gk�l���>�2�{�gdՅ_D��`�@ep�|��֯��Pl��M��� 2+_2�
������C��P̃>��Eă�ao�p� �t��JWQ���Mhj���ȿ���5�����y�_.[q8s����W��GO�DH�)�@$J\��n�a����t͟9��f�ڮc%B�K{~Q@mp<�3�'��
0����E��:��� �X�t���
�����m�&N3��!�U�	[:��z�K��� ����	"�kE��b���q_5<э8�a���w2%r��`M�3��7&�(!X����⩜#b�.Eǽ	�ZnrB�\A����i�f��x��
�P�@�L�� �AJ%�G���ɗ,��m�/�b,h�ae��&}��v�:L�>�'-����ɱ�j�J$����
F�4��	Ib�. :����#����� �4��o�>���u����G�_F��V�	��T�9��ݹy\!9��v����\u���H��PF1��V5�xf�m�Ii݇%�o�]+,A�t|m����Ʌ�Iy%�RE�;�%`bޠv�r�ҶKav�O������a�"��[�\n,�!���vW�Ӝ]��JtE���q��K�c���S�+ar[Vt_~��e�1��(��S�l99��z�3.��ndOM����4A�ͣ��R|>9�S�{�-F8C������^~T�'n�P� �ѡ�����v���9���~ �U�x��pQ����ffȋ�(H�_�r\�<[�%�]�ƊZ�������"4#J�Du+�_9�k����N��Em8�ꮱe����S��/x\V���t�N�B�eU|�ص@W:��*���[:�t,	��V�b�a�0�j�@�Kˣ�/j_�w.�J�v�]���h�'��6���鰀?�����g�6��w6%����� ����Or�u=�qn����ᛋV����%xE�QS��#ûԃaפ�J��7�\�0I��zLx2G��k�SO&�́��Hڈ;PO���x�&d߁߃0�;J��B������z#�|̚-�x�Eq�6K�:�1����S�p)�;�XT�w���en �Jf��O$�Ùn����x� ���e9]��s�:^��{��!H9}���[��%�}�&7�n�\Oj������],,&Y���?���#��B(���pd�$���ic���Y�TNэ[g!�ؕ�4�25�##J��&%�.z�6y!Ҧ������=��W4��[	��� 8}W���J�#:�!GN8��(M��!��'O)�E�G��_�H*a�g����_pv��KU�)Ͱ�1'6��:;Wop�D>��;�����H����Q�a=���M��;Nj��VJ`���f�Q�8��a)g�20qM!nh'����}幑^eq���P̕��K�8j+ ��C-L�����L��oj�_`�:�}��)�Y�R�Eu ���=���V�̚TM��&aޯ�!.6C�� �Q?>�L�v2��fs�+�р��΄�l���b|�Đ��i2|����m&�F��&;�"EV<����t�hgbp2���L����;����[�H���hV7$8I�p~IX���1ti&��>����p�������+c��6�w{d���J�!��N�1�hT:i���6�hD�������b�9��ٰe׍�"[�������Q�J�f���������MD���񚭼���a~g�T���/�y<T���j�M�l��l9��?�s�U���q*�3֤�7ƜG����Hw�e�L"���un8�UBUj����A��9��J���T��\c���P<Hf�O��)����g����sbA[	"�χ�\0�$+�~��� @��#�v�z!<�(��a��5�֛��|����k������IOs/P���*7�0m5�|hȯbh��8:��>W�$��D �7ė�$�ͺ����lȇ]2	�L������݉�Ɉlr�����G����Xh�Т)g�<R��c��H'�{��Z����:3*\(� I1xq�C�2�H�;�����L u��_n�uoJ\W���0+
��oȫ�Vv��h�+�NF&�$��n1Z�@��0�зl6\& ָ�T��E�O��T�K�3�P���Be]T��T(�n<2� S�L]����,C;�8�����o��d~!�Ϫ=(���T�m���g&5�}	K��7�n*��RyZ��\��������gˆ�>8��2�8x�җ��㨫~]�t��`�EY���q�Z?�AQ�D���K'R'�������K�lo�Űe_E��^�z%�˃��U�8�;H�~�njy��j*mhd�����<o�i���UN,�q.�7�b\�g�Ő`�y�X�dغ1���6��I�hJE�dst�Ysg�V���X���va��ޟ&%}u3Q�B;l`�4��z��dv��_9��D��O��?�~l<>���K����iM�X��"W5rZ��b��}hq{hh��k\��pNFD�P���$hgo��wV��*����g	�~7�W�H�yE���O�f���0��-,ƼȌzo�l��q��a|�$Y:h��( �_{���'�d��J��#��P��6Y�Y*A�x�&b63��Y�H�����|<��Ai�E9�E	��FlL#�ҫ�We��Y�q��kna��vS�H��6q�)�w�.�2w����˂���p�N�}r����CX�zȵz0gm1'_M��U�h�F9 ���(��f��e��m�7�~�tTL���2cB���%F��JW�~��}8"_S(4�r��ڬRY��<�-�{�aB|��&:f}3����Hӹ��������R������˧��VC]|�����ӳ��L��w�N�Cbv���ؒ��Qz���v����@ ~aRn��/�~�=�n�o�p3Ym��%W�s���;QabL?Mtۻ��b��uG�8o���^8l
�T#����r7�oQ'���`�آf��V����rԔ�u�;�Y�Is���a\��^��Ա*��SM���>f�1b�����n�I�\��b�8U����;K�øc8��s<<���]HY)�8(ɛ��Eu�${n������dD�����UI��cV�ZWt�~O�Κ�>�s�h�+*H�M�cv^�k%̸����B�7c>C���u0��}~�7��}�<[���^5~�OYsvd�l
Er��@L�[FS�����.r��������N����Ś?}>�6O�r�hܜd(l�`�v�e�!��W3O/��j�B��T����9jd�˪�.bG�C�;��
4�\f9������El`����9�����2�#1z$���w���SG�m�]-�u�p����p+�_K1
���f�2����QW���-f��3xT��q�$��i!��� �{��$�Y\���ل���?*t@R��U�HY'K�I�H�~�;�98_�8�Ɛ�n]m5o�#X���
�Y���ɭ}�>��7y�)����e��U� ��]<gBˀZ�N�L��)��̑��$Uv��M�����i�����!hS��H�,���qO�]q$�����7��C5_.i=C���|�ei%�R���õ:���ʳ|@�%aa1��G�}w��AQ���]s�]o�u7�C�A�B$�w�+�<ܝ�2�z>a��z��#��E.o4�It��KP+����8f�ڭ������u4����[�_z�h�������N�ab��ԭL�1�'ʾ3J���!�t$���������,i��q������P�	M'�̖��󀄮%Jխ�Zy�z�6	jD�%@���8��[��]��+t���H������w3�\m�u�姕`�z.��(�tL[s�tj�o<:x�O����B�/2A7�
^ף�1l���v�9q��,o)U@ ��a��/?�C��B�j4�/�R�k�Ŵ�	�uS�~���@��xLv��Cqn�����w�0��V���Y��s�|���C����9F؞(�0�#r�LZq�'l��6�������������l��EP,��<Z^w�ҸTZJ����)Iz�U�W��B�2YXNNEl�pc����G)rp���� D����/:�tk��`��_a�PDM�tu���b��g ��Z>��V��V�t��b�Pqc��D"��PS}��������=Qb�-%Xw��~-��Is�5@2�ڨ�krZ�����ú.>�l�"v(�Mxy�����(�8]r m$+5�S�N�Ɓ���I������z~k]�W�4h�����B���iD�t`O�{3 m�jx�v�P�o���E���m�'���F9/���?�Ir��ڥ�n"Binb.�47�Å+�&�خC��p_����9J�7b���K.1�z���ډ���b�� ,-�$�����q��mߨ
�� �rp�x�_�K[G/�|��*p��Y�G/=*��l"��������Ԃ��bйic��j��>���EiťZhju_��We���yܫ\��^g��0��'�T{>�e���	(%ǧ��BS�!E�Ï�1Ɉecs,à�>��n��n<�m��M�?�޹O�!�r�k1���5�>3E�M�x�*aR���,&.Y{���"<3����.>x1g����&dJ��v�F��8|�[9񹞿m4���!��Zٽ n��]{3w,>V:��e}�u-EH���M!Qmd���1,�EM��[�D�n�*&_�Lzu�|Ŝ�M�J7l�Ѩ	�E��Id��K�]��\1ʧp �?����oa(U�B��݇kl2�暹�s���>�e�����8y��_� ��`����ݞ�"������;�2L_ނ,�\��d��Cn:�y��3m�B�݃�vrد��Ci�(�}�iQ�a]���~XZ	�B��V��+$>�+��х�vP��T�h/�2y6��yO���	H��"B��/]S�'�$�,���c�g�k�'�=����k������	�X��;�|Ys��RB3�_E��@��bΕ'S�6���q�,�|�g'��u�ʦ��49�H)��"��u�P=������ڑ!���&D/��E@�z�%O��-�
),���?��Bs;��32:�- �\!�p��ak���*>��\��-�g��G�N�g`?�}����J�-$+R�c�����`;�_3`��+�����`���d�=5M�Mk��7�fQm��X
�T:��A�������;�1�G�S��ݪS컿<��ad��V��s%V6�3��$�X'؇����ǡ۔�G}V}�"c"�MB`�WjWN5��qJہ��Sh��m���B�^�¹����$��G���S��V��=/F�Q9f�=��tH;��1��:�r�Ͻ �u���k����9���y��I���JF,T$-P*W{&Ƕ|]$����m��+m�j�sf4�p�͠���G��oN��
��o����w��r:�ވq
R�������f�s���{�I'�ۙ�P���L�foɔ���'�5�)���G�������3��&|-d1�w��b��L)�:��J@VG�V�P��]�����Y�}�#��p�!S �p��z�.�a{��#86Ŏ�ڇܦoC[}q��l�*��Y�A,���u��H�x�T�����l=��������_�=}�U�x�2�s.*�}b-���	2$��u�ۢ��w���݊brQA�d��a	l�ڣ���$_���k�gCb�#�R�N�۹�QA�ߝF�^/��sq%�E	�ʜ�2K��9��O�`-����o��6���[�dv��<����2g&����׋�z����.0<�=�2��z9��u�vJ�'�K8y�"�T٭HiXYC�<��q��\���u����߰��H�}��}�rX��^ÊV
(�e:��4l����ˆJq�::I��C�R�z��
�M�k?�ܩ�>�F|F����0��uTkM�x�ߒ�<1M�B�?F.�ev��m��J�H+*������IO�vѫ����3���@��iKU�g��y�}`���_;�qR[e�^�����s2�+2�����2��G�t���A6w-��K���?�rG�ca�ѓ�2��ܱeA���o!v���m��G��V簂��Xt��d�F��Gtg���'6� _6�⹳�n��}W���f-Z�}_�<\�K������oح�e(Fl�\8Q�u{��U{AD�g�qs�+w��G��d���T�|�͆�t<�O
��L4���S��M_f�C�T�38}���5����7YTB��KQ+�9Ȅ����@��
�P΋�L
Q���?�ѨP6��h�7��śf��x��%9
�K;��6$k���E˷�������(��^|oq�Zץ�A�w�9Ɏ��K��zԣ���������"u�z��tګ���wZN�c�%�M���J�J���T"F?�/���U��̒	�J�|���ŀ+7T���M���z�EzX71�!J���w�4�_��#�������uMpZ�v���=��aFd�� ���L���_�^+Z�jP��G�C�R�q��Xu*n� ��aU���O5G��R���G�r+@33x���ˠ���OAh$�U�؆��ׂ��2��a�
���f�g"�&�Y��<$�_B/��#��~""8^!/��{��0_X��� s�w\��nw��0n��O �����1�1l2�h�����ldF��Og���7�i�a���o�]-01i�L�U�)��s/�h�J�};�[^=�Ii�	#[vu#QRa����w<lY���2�������V�
%��F�u�r�~�a���j�V_���
�D���d�\�X2 ��Y���yV��H��5j�!�b�]��+����?�	�#;E4��iB4�r􆇓�iM���=�8Bb2cR\py�޾�}�i�����o��F��a�[�^A��B"�������֓E!���X�����ֆ�&z�#� �L���\,�,�Ly�s��S��'���1�[�l�������rb�倍�����,��V]�ţ�v<�ב��D�RpY\厣����y�,s?>%�3����P@V�N5>+3U��=�=���Z� r��^�����[ҧ�G����0W?u�\޻��t1,�V8(���xۊ�����G�܈���ҩ��v���o!�[���~]�1�'��_�jh�ֹH��u�:�m�^�/ zʆ,�H��kse�80Q�j���yMO���xW�ǴЅ�r.BW���2Vsr��amъjTq���ѱb���#��� aP��χ�f��]��)�ȵ���C�c$)ƫ<�%꬜(V�>u^�z���7���� ��A��^伳)q�B-޳���%ݨ���R����K�������B�!�Pr���ګn>�*�	�e͐_�s�G��5�1�3�rl
�f/�h��޺#'�9�C����#�Yqo֜%��7�����`�m*�Fnk8li�1��DJH֩�ܴH�)�� f���m>�&�7?��)zUҕG�(뱃䢨qs�4o�,k~������&.rJ%�hδ��'0=*�S�:'��T�aF��UMv���j?�����e�A��9�H"�!�	�r��PO���o��N'�]ߛoN�a�Rgyp~�6�$z�#�"�.{*�&�7��r�tev��|HG��̿��Ϋ������v�Fѕڳ�L� 8�m�㍫ ����o�
��ӿ��W���x�,Y��L�p��P�$|��1�2{��y�xU�'�^z%Y�_��Z1A͗��w�M��X���� 0�����2(?�j����kyǣL�~Z,���v�@�Mg�J��t�7�i�sT �`���x=�j�ڰ��w+f��
s�)��xQ�G�aF�G̼N	���'�3�t�^����´@ӻb/����2���	3T�#�������jG�2Va�Ck�St6s7{J��cn%B���@��6���|�QI /�{�$ )�&�v S���d���A߳��ߖ����2v(o���ƒ�Б��Q{N)��ypW�z�I[M��������.y�~A��~A�S�u�3 GY��nLM�!���v�v�B�W3+9�Y�Y�â.m[��0}���)}�(��F�.��Jeh�3�(��Ҵe�i������G;Z����\E��*��Sc5�geK/n1xI3�X����Jչme�T��@��~�7�<��,�З3�}w�"��p�r�G��e�7hj�UkL^Skgyӏ�z���4��8����X�PO�i�0v���9�����yrD�u�p^�-�nG�Ө�rw��j��D�О�)���rBGvT�-�	}�EY�,�N���`?��+C
缨��qv�@��p]߿hW/҆��A�oq<�������QIOfO�d�&��ҧ*�rDJ��XT�����J}�F|�p����͓KE���f��h(xP�w�$F4;���̤��g�?��,�!����{��S����a~NX*�[��q���/>�����lj��8����)H��PK��ŵ�E��P_�����,��?q�-��s�Č%�j�1����7Q�UèE=�Ҙ�x��&�p6��"oM�Fe�5*Ê��*"!8*Sv��}�A���X;CWI'D#82��?I�G]y`�D
��6��C0��%���xm�o%�7ҝs��E?��`��"&گ��ٕ��qv�/�pqa��QS�$��Bd���I��\g\'�`JJ����n<I{�x�GWU�hp]ӈv �Fav̊I�-�}�I�_^��:���B� ���3�V_'dNaC�:ܽ!yS��Ѱ8P���H�g��������W�E�]��"��80������o�v@8]1�I�H9:�Tlqi9�[�Cw��d,7P�7�3A^u�5P��\�Ϙ*I���h�Ԫ4��s�*�c3�@m�����>Ѳ�y��$��p�*�����q��fgp���:�$^o�@��常��`ɵ��?�KZ	8��Uh[����jFI�?dv>K�;��|�� Ӿ�P�=1��ܞ�D4?��b�PL�ȊgEs�2�Q���+	�W�����Mh�\��pL�-�o�;D���§8 An�x�,���?ɩ�N��	��Z�C���?�;%�Zۤ�淴Ԩr�o����"�brV%�,�~���F�����0ot�A۶P�?�۴ϙ�4ce�����eoC+?�,��2C@�i-�fp��.S��,�űB-�o���8��2 bSө�Z��;k�E�g�����T�fa� ����~�h�v��#ݼa�;�3���)<#�;O�;�'�	�U��<����N����Rֶ��+!�� �:tT%�9�Q]a�K�$���&���� 
��3��z���_-e ���bz����п���'y��U�B���@Jfp�{�ѻ��5!$�-IP�i*#�%I�Q�)���wh],�%�R�'(�9h����gF��`<cw3����&)ҶJ�0�m�|�`AR�ֺQ(��9*�K5`��}���9����`C��ջ�iKl[q� >�X��,��Q��ҷn�`c'�z��@�s�qJ_q�@=J�.m�0F��\���=������<xG6�tĐ%Q�o�`~���Og�`��a�%C�Q���-��(e@���Or(@ҳH=��
�����\UBN/��v�%*��ؠ9�t�;6{[5*|��3�rΛg�@�9�G�ع�t �
G*��.�K`i.L#�`�Qt�j)���s��3���K+�<�|�ea�,Y ��Yx9��|<�*ѓ��t�Y턠���Di64,R3���hQt�
\�Y3|�ϝ)WԃC�l0�ҿ۴#;OQ!{�fޝ���a�Eۭ��ќ5�\��Gq�۔X�Und��Ib�@�Z�����9b4������:ݨߐ�D�;=l����!��$Z�/�	�P��6 왔����Vk] ����$2~N��	��4�>ǰL}�+�����Z�%Z&�6��9$�g4J�dK-c��=u����a6p)R�L�
UC��
l=r�d���MXzK�/`Nb9����R���ρE��(`'M�kQ���/���p�P��X	d�I�s�\d|��̜���2F<g>!��&Δ���U��p�K�E�U�FPx����b�Us[4�K�`��rF0���<o�lp���ex}�t�l+���նGT;��9K�7�?Nn:+J}���Z�c-a�s<�a�|K������L	�n"T��� �o���#�*���i֘{���o�[�-�_\�y�{�m�T���w�� lURF��YkHO��R�&�1�0�Aj�uf@�"vR{���	�d�X����GU� �r���"��Ա�jQ�-v�6d�����ۚ�UB&3T�YD�qx��TH�^��R��
$p	n�E�(����������_7���Xg$���_���hD}��!�[�A�I�D��]�/ƢFR��؄��L��@.;cq� �t�N���Q�"�M�[�(0�	�O-6�P�/|y���V��'�zF�<�7v ����5��ޡB=�$�X�@Z�\mEE)+٩��H��Gl�z�0o��X�}�ҢBn��z6vA� a�ec�M���+g�ҏs<� ����.�����雦9�}��U���\FZ�	^a�fJZ��g'鳦�}����~�=�C@/7^��cQ�B��,y��ڶM"��5'�S���Ѐ^���>��.&	�������m�HȦ��U�z�o��<#(_dS�̜G�+�#�<��3�Z1���7)y�[�thQ�^�����A3P��.t�*ݱ)�� �R���(x�)NQ�֘�DX�w�\�D�+�f~HP�a���FJa{.�����w���e�g�[�'�,�R����J�&hT��7P�k��ޕj�Q����_���RU��� �����!(1Fk2��9