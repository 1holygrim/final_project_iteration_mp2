XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ܦFDՆ�c�<�x�Kƅd�3G���c���_ �غ�[}bWs��N��P�a[�AT^��M�l�$�s1�L�'�eL ���+�"�����������n8����ӿ��;>~3�܏5��Y���X;P��&f�=	��=��P�[��9i����B�<��e�ȶ�i۹�0��3\�
��\�c;�c- ;�z%`������4����Y
�2�w"��J�I�͘�r�O�3�N�i���A�߯ύ��+Ի l1�oƂ�\z{�2�7��=[7�KZ8.+�L��/�9t1=�Gp�Q.��k�{� �ʻ¸�M�1T� V�Bj�K��T�S�:ف�����M�kvMl�	����s�Cu�h"��Z[���̕���V|�L������㯈�e>e��Xs.�%@�5S}���r�Şf��R�7��}:Ȧ=���J ��t�Fͳ�(T�d�{�ċ$�7N
��Ω_q���=Kvo7�W9nN�h|/��
>{^�\�!����a�l v����F�:�?�9B����Lo�ah-T��2qp��wOAQ�V��W+ˠRlvf��6~�]�d�:���Y{I�=��(84B���ny��(��q��쫯���]W�"Hl�8��Fǿ:�C����U���	~:�^�5N��ͼi�WXj�~i)�0W.V
+Ё��A�SJa7ջ���Qe^����\�������tV����?\���f�NLJ^��o����Ц���@�m��'\#V�Ŋ}����w�:v7!�a�f<b]�XlxVHYEB    266e     ad0��0^�%h�H����4:,ōi$��0e?�"�P���0@(nb��k�aĴc�0��x@�.�t��$�2!��w�[����a:�Řn�5__�C�aZ6˴�v; �.�,r�vύ����9�ƣ��]3���3*�D:�f���˛��k�����jу�1��V��8}|�[|���y{IV��*G�;����m�a%����;Y[�EΝ�V����.h~� �Y�Zn���n}�;xY[�"�ku��~��g��@�h��©��:�ի�\�
�/�3x�=`��a|F{�X�����և�,)G[~�8.a�,���)��m��|b����t@����u��$)����4w#vF8��^�])]��Ҷ�����\�1��p|�2�$�NV��`�`��ir����'VF�b�WfsD/W�Y6#aI?7+2o6�dA/�Uv�s{�g� �D���q�� �Y���k�j���R���t'����`�җuR���Û��� �������L���:�B�@3L\�lWe�*��s��=�k�]�������Ɋ�B�YV���©")�1=�ek�I{_�\[��>|�"#�]j%�-�~��թH�Ȥ:G��,$ӆ��HV]/�i�mC�Au��׹H�c�u�W!j%�Ғ�|�V1',�OO���Hj�eLf�Z�}4�2x�$C�?UF�0VP36����o�Z`�[�n��L�8J�0������[��H�pb�=HN/� _!<�*EGt�9W=k����]ۂ�!z��41�ERa�dr��WC*'P��1I���u���ɰ�%�w��x�;ʞ�|��΄7����j
�BC!�R^)�M���*MT��`���g�� �N�~x��E*��|�,�b6=#��P��Y��:���]�䐤pE��pE�e,%�$k�I�r�`9&�,
�N�l��H���&�Y%���cP�ax!�zDj��n�v�4���#4ȩ?]e!t9b�E�SQ�[]o������9��eLl�|���^
��c6,`�tr��aV��F�{�%Ku��"n�;����`f�3�A
�w�|�����_�N!d�:
��yt�����:��X���� ���܉����Z j8M*�Q�<L���C���4e�f�1n���C�I�/N)b�$��2������0y��r�]}p�ћ��\6	�-��� /20�{Z'��۷��>�Iz�ՄZ�����>�A��Qn�ָ����6���0���Go@���i~��"w9DD��Ղ �$@v�|�*ȉ��r���YB2��T1��>���U?[D��^I�mqp,�����iE'Xga���2���'�u�ɓ��C���jJ�|'��Ӡi`� �e~	li�n�S'���ug��5�	n�3��}�aɣ��|S�6��z섲p��*�F��y�:u=M��m�|�
�
�y�@0�&��	��T��ȶ��JPҊ��V�m�+�P�I[e���Y-��cd^�	mw���yUnM�j�����%��~>����N��CV��A���m��!<^�����X	��T�y���܄dĀ�L�Nl�)���k�U]A��p�uY�=C�����R��ܿ��\՗�ԫ��|�)�\�l%/�<�$r�r=�F����S��;��Z����M�r�H�э��;�ނ0[[%۬�}��e�����-r`\��^�":꘹��YQq��Y�uV��Q3�@I�ݖ}{:�R����΁,}�K�)�d�#������C���c�s���ca��y���G��4��-�쭜%�,g��>0�ϵֳ��Owݕ�����B�i>����|��K��d�-mZvςg ��:��C�O��n�p���Y �p�1�����Ȓ���es({���--K�L~���t�}4�����-�U��'�P�dZ5h�O���?T9�C�4�!�E�������N�
jY�,	Vu�D�]w6e�GR�,l@(�V }؅Xp2����Oci���B� D�e��`�>-��8$Ђ�}+�Ħ��>`B����\���+#�*���F��,R�Ə��Ѿr�u%ז���8�3.]�B�GVZI���*���ds��e����:��Xp�#^��1 ��L�ǖ6�~{'�v(8����fn��: ��lj��tYdơ��|?��Ӻ�qՌ����e	l?S�h� �5l�:@%�Pu	�/)T��� �S;�i3���(BÙ��{\������I�j���9YC���^�D��c�vR&���n
�$���|�y �>�mh������$d�����?>����3tF-R��J���l������I�jC4X�Y���d�J�Q�2�'F�$�U�dz��
⭕����
\�>oE��N T�1毞 ��"�6�����&��n����W��b-���iW��$��9�2yo��.Rk�#2�i�VJ\6Z��l��wXD���IA�L�i�%x˾ˌwa�Uճ��iV�OV���Ad���8�_4�73W1?fjhs�V��O��Bt�1����t��ē6�E��u�@` �2�߳I	T��$q��&�7����*��<�^��áVH��tR��;��C����K����b�VN��4��#y��u�����י��~p@�f�M��0�p��ڜ_S��sG0O1�~��S:}�P��
;�~����C`�7*��;��G"�mSZp[�CS[�3���_2+�2�z�O�/����m����̢p_