XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:z}�+&?q<�W_2��N���c�0o��7�:"�`�pξ�� |w��.&_��V�0k�;��r�^���N��p�����\��٬:7�A"iA�;U�B��Ϩ�������b����֟?*~����Sn�����p��Ї��#��?Z�Xo�l:�����MQn�lGls��p�H.����f"�Io���pgo�bj	pi��6��~P�#J�)�m�� ��;^�y�)�ZLy{�5'�,r�_���� xo*�J�E"g��3����G=e��8�.XJ�K��.U�@�b��|�Fw�u��%��M��t}Sr
=+!Уi��c�$ll��.Ӑ�����T��7(*�E}�Y��Z���+m�8lU�����W��N�V���;b[�řm���*��s�&���9���^Y�u���+@J�a�Ƶ����r�.���̝���6<���VW���4�,J��9T��곴�悋b.��k�#/-^�>Vo�kCOؑ��)J����bG'���E��j=�fC�!�!,���Ԣ�ay�ĈdE�,� ��E�9}V������K�����HS�R�d|��p����9S���Q��ԫ��eg`����)��M��|��/d�%2'���!b��4ޅS��l�����\A��!��s`E�[&Cq�9R��TRnT-�Q6��IO��~�y˗�*FÂ]�����a;\ڂ�'��2����-Y�x8%b�0�\� (� �.�|�F��|XlxVHYEB    9852    1d10`K�8�Q�U������o�2@ᝧ�6%�;�U~����:H�1ZZ��c�p'�ݕQ����Vu��i��"<�{�gI�.jU�6��H�.6�O���B@k]n[��C
UG�1eX�eA��D�B�e�AG�D9� ���C����l��<V��M�?LQr�s+�ǉ:�G��N�<�5)]�	bLj-��dJN�P�o��:{u >��{#��h�u\���K
��uP�~ah�Lf��sҨ)}���]�Uh��K�C��уƽ�����^������hSQmB޴I�eSV�;`�����U8:\�q��ݖ��6��`�|QRX�mim�_�uH���T��"�3b�!j"�
F���RP����g�4��"����_�6��Nh�ޙutGGR��8uG_�+�S}d{d_����8ZM��"Y|�����,�Sx>�-E�u"��b�D�2��@^������o����T
��`�/5��3�s3���ӂ��|UC<~�<�x�i��D¶��:���o�����yI��>#\�,7H+8X�H�S��t��5�51N�b�#���:�ۋ]��*��hdp۞1���)8pv=�ܬ�;� i� �уXu�dxt��i#��m����x��I�s�G����I��X�l#�Q�q�^�>����5^����	_���e��e[��8�;���O`���A��ޱ��_]R}r�/�׋���]:�f=��Uq�����c~Vn(CD�`�xc.���'�& �K~f�������2����������Y,�Tay�E*K��a�aS�3$vxPի�޽m���Q�N5˰� �ܽ�J�L!c.�����r���Ct1+����;a	�˖Hуa���M|CC��@�g��(��8p����4:�2���]�䊲i�J��(2�Y%͜g�2�{oԑl��|U0��`tz��%�&~���Oy��C"�kz�rl;�(D��:6�e{�(�ڽ�$�l��y�D��ѿ)/@�2H	��|�Ҋ{�hI�7��TbK^W�����lE��o��6�Sރ5��5�iD�`����|�a����I�"d����T��.��J�Y	����ZM�� c)5�6t ��G�u(�:3������6�����Gwݷ����Z��&������!��S -��f��H��(��j�zv�qz�A����S���x�Og�N����X�L�.��h��͛��IT�-M"�N�,r�l(�����q��K�dB�Ie�U1�A��t�д�cC>��jA�eKvM.�z�D������H�w�8�Ԏ��@7���q�Zn&�E^q�|V<������ ��5��P�����D����]������i!	(T�#C��ϲ3?�R�(�W��O�#�?+82kr��*�O�E�@;$& ��AT��N���׭��*@�]e1�x�asdRW-g��O�ƶ�<j����5:$��������o���5�I�ܞ���]�@A�� e��{�
y�om|f!�G�ߤv�jI�.U��y@"[�5�.���[~ B��S�N��B��j��o��>�.��x�͑l���8��ߔ���h��qQb�P�5sְo���c��<�����(�� n�§���]#7��F���]��
>5��������'Q5�=A��'ZS����yύ��ǇxK{��l�a��z�M���J�?' � ���sKYܐ-��|0k4���~�}���D��\��zws|c�ԌL���sa9�&���g)K>�Q"Ӿ�+$�H�/]�j�M��Dt߇���š-����L�\�m��jv�'6�c�S0�F�^[���4¹�XJ�U�(]��,�SH��$ �!�A��/U��S�d�l��� �&0��[8	nr2���:.rT��3���9�Ș�$�Sn�y?��x�,H��EFcҩQ����,�ݶ�X!�G$���?#Z�k�`��O=��x.�HMw�x�K�0#i���t���F��_�Υ>��R] �}R	�����G��Ui��ѩ>G�r�ZZ�B��^�T�x��m����m��|�´���:�+đ���,}.W��� n؆�[���ױO)�A�Z�(׹�+�B��oT=�Y0~�р�a��P�-��(��27sڍC:�7�N2���j*患r����	$*K��%5O�w]�Ð?k۰���_9�:��3�ח�d����h�Fӝč^T/�/�lX�S����ԫ�0�=U�r9������G��;��z4���R���g���s��E-�uֆ���sd�aEpV����1�����9i��1���F"�FI͏4�J�A���)Җy��i�-BT8.I��aR��(�S��T@6�T,�'�Ա!+��Ec)�u$^�����6���Ȉ�=���rcr�=���sdnn��X��E��Wȧ���ԃ�����5g�~l���KN�
��xD��ǆ���dC��|]�˷dy�N��ؾ�s*AO�O�1
���L0vt徠&��q�t�����r�^+ g�oԮ�L,H�g���[��ͧHǭ�Pj|�}m�Z���X^��X���X�=nٗ\NqW3�e ���5���8r,v]�7�O���L�#�9�vK���� �T�%s-?o3Ѽ��x���m�Š�Tw,�P���� �ѤCO�3Z�'��
��T������s�Y�8�;}�>�����*����ߑ�,��;d=zݝݒ���W�$2��V4;��Ǆ'�1���=Ǯu0=h�-���h��IKQ����\��X���p6kk/_�d���=�H@0&���Wq���\yX=�lU��t1���g&+�,r��M����\#mX�;f��2H�'����/7,�͵x��ƹ������շ��Z��`,��C������j�z�i����������	��m6��t�
���� ����g/��Ν}e�JqOe�͚�б��$�wٜ	pC�8`��}1�9�Zp\H8����@�P�}3�Ƞ>:s�t�C�{��k@�yz#?�����:�t��>�������눓gX7y�8Z�&�,�0�EV�W
��Y�6����m��-PEY=yo����{Fȥ��aC� [����Ѿ}u8�V9d4ydx;���HMY��	\���]�9��D�x�)��U3̇,o8>�!�p�y�S�I��vQ�������'S�W���!��;�^�t����c�>QS���hgWÆ`���+#��@_���Q\�XK����v����J ��̀���<)v
Z(�к�@� �G	�{'��WBIq����*����*���y���D�d��"5o������#�9���o���oe��&�9l�U�;�[��>d��i��)��u����pھ�2@��5"�<�F�?
n=�K�o���4d]���z����vUdI@A�,vy�ή+�cmJ6���y	x��e��ȉ����T?!狼'`d�����̷�L�5�é\0����zv�F��Ň=
����+�k�w�L �g`��:�^�|up���lm~�{-����3�'Z��$x�������Ww��7�\�!{�z�M2��^� �XSc�Vj`teؒi%p�w7.JJ1�k�1�++��J�v��m���n���j�)f�_��������;��3q��չ���<՜"c�g_Ł�OK����حm|�2�h�li�� �mxI�۞���<�2%^rE;���v�ĵG�� o�qos� 3I��Dd�L؉��7���or� 9{f��B�&WG���4��bs���X{���uÉ�J�=�6
�m� �ߐp3F����>�z�vB�+�&��CVAt��:IG�{Kź��>���o��#E��UOW�kp"��4�C����4�9��k��h��4R���Y������4Ñ%�jڈ��EL1沬5(���o�nT/��8����[��2���5��A��U��B���߶��d:�B7L\��L�'y����X�k�A�o�h���1I��CTW���*9^�A{��-��hd���^mpT}�vک�,:t���>a*�	J!��̂ a� 0��@��L�W�k�#�Y�L#�c'�����{��S�:�DM`�d�V��vҋ����!�z5m.������&�$����=�������+���g�rC�v�'� XoF~@�B7^���M3N�xA�������@L��	���'�Vp=�͌��/��XFr|�F��߶z��J]��m���<v |Q5���J}��*hދ#կ.�ξ��Ӑ���̡��7#; ��{�Ow���r7��1�F��a���;�<ز�ÃA��u��`���XDF�Ƭ��D�v�\��rl�0�P��ÔZp�ģ�p�S�a��4�7^��A��L����3�ȡ���ӐH���_H��3y�qd�H� �
���H�37|\L�e{�c�^�"V�[&�I[�I,"�skE�>>T��V;�a����q��j�� �E�_��
<:��{[JyYD��A�F���+JL��X?����=�:�sZQʇ#Hq�AG�t�]���� ��2�[C�J�����%���wL@�=�^ZĔ��A�0��-����?�"�O����/c�9��M�1�GCXE�/��ܦ���?6#eD��bW�(P�\G����	�H�����u�Z_��q{Y�S4a�T��_D3���pA*J�+���r'��¡�!a����7{U|/�ٍ₌f>!��M|B�d��O����pZ3�U���=�_��W����&8���(c�>�ޒ�_�Gu~�5�M���XC9�!�vt�q�qsy�6ζ�;�Υ�.4YD��*#��i#�s��$�|D\0��-:<���z[��D�Д�qF<8y����%�R�s��Ki٩� �4Hۼ�9�W�>���!u�DR�z�Ƿ��C�>��IF2:�?]�w~�BA����\sK���j�X��in)piZP�雡|���F�t�qw�ǃ�B�>n����w\�h��H�~�8T�.y�"�Y�Z �[N:�@A��B��#t�.&�I8��梪�V������38wr}���>!@�4�yCr�zS<l������w�Y�tw}=$�'�X˴����F�Wӯ� ȋl��t�U~���s�����-��>WDĐ�v���A�A�H8��P{�m6���_���>?���a���x����h��	ց����v���#�qANC���5�U�����.��י�0��`��M�����Ҹ4e[��p����`�����]�Z~M��;hO��'�-L�e}g��1��m\�D���y��<��aҀ�,��}�j3+�D�$�ߨ��i�a3����32W	T�i�/k�.��+�wl�ڌA@��[�o\�8��|>�tR	4Z��
��W�CȠ&*�C/q���rcSGg����{�.��M�m��-
�R�7g�у�a�,6ЌjW�t~��1�^���H�Rw��Bz/nA)��g���t���m�A$��F�#H����v=��'j�\�%��ʿ8�����SV��ً�9?à��6���dz���s��z���5^�9�L�R��z��fO�wrG�\]9��d��d�&��t;�w~�!3|y���m�b�2 䗼kNݼ+e����H��4{�q&Ό��K���O�a|�Z�-;X�vC�#!�]��ppf5�t��^!W�X���ȥ��Z�e-S��������C��0���������x>뛺p�d�w����,8c>j-{S'jҳ(�)�:'�w�?�ye�r�"�M�mBX�͒��\ag6�2m�|�8� �����z,���p6��H�L��x����#���-!� �l(�ĮB�7���0�`Z���PsQ�֣A���+3B�����w�j~&�c��	�&��<g��FJ�
�`���֠\^�:�t"�OB��m������c  Eɡ�3���i���5�E��xM� �CI}�GZ+��=ت�g�R�䝢B%SVu�c�����S�����oxa-�����w ��ԍ O��/��C��g�Uc"K��!���x�Jx���vL�@xt��Π���<k$����x>FŖ~V@7�v����N$�}�������y��ؖ2Ӂ9ȗ�녁��e3^����Ksl������zbU�NE�А�: ������u.K�|���|�I\��丠J�D;��ml�;0�͜�wԤ)IS/<s�e�/e�Z�%�����Cސ[G*�w���ҝS����0�Ca����%��+~|K>�I���5t� 2����p�K��J��Uwc�Z�:�2Н�::v]��\�	�^�'b�ӿ}�R��M��������x�h����μ/���M`���s~�X��u����7f��]�K'��C����ƿۿ��iԘ�1��aEA���B����ž��~\�'�n�6T�3\�32�e�r ���/�<|={��0�0�����0���2:��wG���j�j/�*�K�>��P�#�0l�7�t�Z�PO����LƓN�����_UIm?B�{O��	%y4��B�t;p@���9�����)i�;�ى/�bۖ_S@?���K�m�
""��_E�7�@��x�#;������Z	��������7��V�|s�����u��*6`�j���Cz��H���L�@xD�s����BϜ1r���:2��l��R�_�Fc��Y�6�Yh����嶇{s�[�I��[��=��կ��BNG��ف�"�������gY���o�L�`ҵ`�њ>&|��E�j6��X&mLO��FAIݝ}ž��ۛҲ����N19r�U���'�|����O��	'��ؤ�v����T�Q	6�}�NBB��&��.m�0]�\k�a�i_�#)~�a�O�@�,� ��b��Zΰ	�����项�H�:|ng�.�:�=,�KP��=z2�v��/����`�j�cb�$�8&J`���Zt��fuW������w���1�z��`�a�[���D�5*�폁��zF�H�PZ���f(��&��񝅃��t�#� o�/�X��J��B�-��whx0�{8ܧ�0�K.�t,`��q) �5��,��bn.V�%C�r�&��@#252`�,Qv�@=�m������%�5����cO���h7P5���1��Q����2M3 ��ŏ:M� g"zX&���2��S�-��O