XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������N0>q��OpN�`�%�a"J��0��������"�J�]B��A��[�S/�m�,fS?5a��5⚕aF;�~V�ڐ5���\.� �$��	������+رv��?6M�$3
��.P��b�p�j�;Ķ�;#5�XmI,�6�-NN-��H�F����n��������*�mvϝ�d�	��&�x�`r�d�^��,��~5%�B��<u����/�n�
MP��1�x
x�1xB��ȣX7Gz��)	ɘ��)>X�Wrb��:op��L�"?vf3[� j�OjK���xЯ_�;�+��ᬣ�؇�1[�����Ѽ��ځ!����-�~���'=�(�XV��}-�?i
0�6*�U�cB�-�����l�v��l(��+]����Ԛ���ϭ%Y/��T�E�,�LTo�VE�����g�C��!Ԟ@�M��=H���fSC(S_9��]-�U&]E�oft}�|3�����,����P5����
7I�0~3Ѡn5Ǜ��6W�����V��A^��1j��IW},zN�;{&�~���B�y���b����?�����W��>@Bh�,� �s�Ϳx+'��Um'KU�U(�U��g���0�J��=�b��K��:�+`�2i,Ϫ��6?{f67�>�&�zMc	>���[%�!<D̉X�e�A'�h��5Y��hlǮ7#�������S$�m�ב���4⤇G�u%x��pO �)6���w��T�^�B��?����k+��$����TN���au�XlxVHYEB    fa00    2840}���mK�[#$��(v�1?�A�x���Q-��S��M��赾�1s�͌{�w~<��=�Fa��\��B�l԰d��������*��)\����"�i�G׀u��	V�|2�Ŗr��А�C��,�4�\����a�
@�Oө��Ipqxw���xX���ONit�'��l��I�ķ{mcN�:(���ʪV;L�A�t�5�hf1�qe���C��������?��S�}m�h�s߅]��/�3��[ C�W�|B���+yd��p0�)��F��/X��feg ~d�-��m btX}�)<;��j��y�(��C�u1�P�����^-���Z@Q!&0����8]R[��Q�f�#��	������ӵ$S)ؙ�X<�S�<�Z=�b ����k��b�}��O�jp ��0Čd�Z�� n����j5�o���CBG}d~S�y�����`p�f	+����q�ͻ����j�%���5��QnL�����[$?�[���%����lg��g�Mg����V��4[]��~c�\n���TA�r���E4M`<��]�"
�
	�>��<��)yr��>y]A��J�=��I�#�,q|����o�cہdUg�EU��>&v<�=$�ׄc��߁"�&a����`��ύ���!o�&�/�
8����n�Fę>�	L9��8��FN^�+�(�}O�)����U#F�(��=K�4-6FX�*�N�,����	m3=��ph�SD|=�҂�k'�Ӷ�6 L0���_
�`j�Ry;(t~�����V��]�(N��"�f��H����~f���Ѹ�a[S�^�a�O�֒	C��4�lY�f��2�5Æ_�`͘�5��Q���m��@g;��"��R�b�cH� ~�E>u[T�'�&t)��g,Z���Dy"=P��!��v��7�>�z��f������.X�:{�(�]r�I�����N{`��,�2[*8u�T�<� �,�ۭ#��������-	� S����)�C���Uݽ^%���"� �-��p��}�G�����2��Q:M`��iy&�!v�Ϲ��Z��!�j˒�k����!��`g'l�.H���,���ƈL1t9�}<Y�qA��͢;kP+nz�N�%�sTt���Ȇ�]�v4���oH���o�a����lO	7�NoC���?mvv۠��dĦ]��P�O-jR@w��$mENΕ&��i@D�-�'��Һrg���`���Գ�2̨Ss�>��l���0�������f��^��e��.T�5�"NN�ߌ�ذ�Z·>�yM��&��A�`�<bp+¤�u�V��=$�QZ��x1��IR:�<*�gx~p���ځ��lt�耪;�P���*!������׶��bo�P҅(f����	P�ao��L���p�L���?�5�X(&��?
sK�54�Zpg;Ů��Y*)�1�eKa:�X����}$M�7�jh[fިz`�oZA��>�iv"?��7]��(��Ͽ��F�O�ALa�J�����XP��s%��>�<�t/x��d(�rf��o�e�F%�5d�ǂ���H�͉��Z!���\���G(�E�r�m��{����`��B�2:�_m�6��:b@�|c�&���*�	���������$A���ԡ���ð�P�k�#��`t*_��YTd䗸�Y�"��I����2�Z����B����3Җ��}>hn-k���b��lP�{gd�(i/A��cO�VA��Ö6sf�ZI���̽�
�O3J&�X�Z����¡"z�֠���J�>��d�Z8'���S���	�1�	�=`�
4�
Yޜ���GN]El���2e��o���L���]��}t=*6�޳�����WxY*ë7F��*�{�_#"7��
;�B�_D�A���%]@���Ɍl�C6�^��
�>����wO��K�
��vw�$}�I,��-<���aNY��O��2i{���k
~P���W/CZR5�+�NT1�.쬀��S�p݊ǁ#tq<Ï=p����"7,��B;UB+�ؕ�y��_HR\خ�ې����>B��?�~��m~v_�Y�Ö�VXs�8��1m��T1��t-1]�;��A#�,�6��H��>_f{����-�����ZT`�Ɗa|����E�Ŗ-)	Y1e;�]�����[�M�A�u���P�ӾR�NEj�JwAb���@듢�O~����A?l��oh��o��7AA)Q|�uh��	������B$U}���}}��.c���,�٬���I�ńl:��m8�)��]�H_� �Yg���mI8�/\�Y�lrR�u
���Hq�o��ܤg��˻=
�Mu��I5>��|u�.�"5�B�3@'�M���2�hI��I���	��,�2�i0��o���z�BI���_���b\HL�'e������nÆ��,R��Јt��{qSpiĤ�-�@�;���R:}꟣��Z+���;f� �-O���&.X�(?򋄓Jo�$I�9�9 f�hX����j�e�N�,:?n��M���ٚb#�5O���k_�&���w�e��.�\�"�dDɴ�Ui�z{����5r2[!�0�Z�ȮV�#j���˺�X#4����I�7�EJN�|X�g(����Y��o��)1��}��%�癝�M��o�vz	>�M%�JS�H%i�K�U�)+�����DӪy���A�G	�24�Q��(�Ѝy��r���a�u*]yzrV��k�L�k-u���XƱ�69A��T��
����[��؅w	����i^:*Q�zx����*l�0{ �S��#F_�d��f���x�N@��`��sV1���oW�@lbí�\�9
��A��[:��գ�V��E��A�K���{�t��
�x g����.\��F���`}7��b_n��6�9w�hz�l���*�����0.����Q��#ĴB.5�:�s�
٠�AeF_Zϕ.ر"�%ͽ� ���\K]�Z���s��V���lTw�G����B?�Kh��I��W�\��/�O[sd\-�N-�sw��{7M�e�I����y��E�-w�f����ޗ ���ZO1�߽�}��s��.��7�Q��)D0����"/X|�P�_�8a-�ݠr(j�bP�H��ڥ��>�;:�}��,�$|�@��E���ֶ��46�wCq��Ҫ�v��^vk$���у{qzGBB�H��uu���>rW�Kw������i9l��:�L�u�(�<O?�)~�e˕���5CX����.���.x0ڪug���J����:^�)nJA�n؁6������"��!`+��C�Y��.��,���8��8��خV�]��Wt,�R��g��ɣ���v*j%��@�����8aF(c �k�/j�8 �y�2H�eZ��
�#�p���ST�1�BuJ?-��:.����Hk�l�眆��\ik�h�ĥ��q[�w�Y�2b���"צ<���f��������V�a<�V��\I|$6�g\\N�e�j����Z/��.�rY0��C��ZL����S:T�D��8�F*���ߺa}�;�ܯ��)��|+w�������y�ߤ!�4���"�P��8duu�y"7��ND�K#�vE���6Vߎ�����E���MkV��^,�(���L�f�NR�8�c�=�UX2ox����ku�C��{��3�Զ0��h�)��B�\r숮�����yb��<BI5j~�}��ׯ[����ww�9��^��$�s��xƮ�AȨfG�8a��K��.�'�љ�[�Z�@|�����Ė�������� �q5��<�Ϙ�U�?����}����dq���5��($�g�CoQZ;�=�7��z�X���@.�%"d��1��{��%eTTQ���*�#���g{Y�VE���v�Mn�C{܏����4f���C@�K?o����!�@E6��T�۵�U(�`�G�W���'�N���#�����%�����i����n�*��E�|=�"�j�r�ǁ��`���rg�P�#��jI�ʇ4���\h����)3�=y�i��5AH�[1^�2�*��(�sSN�ɴ�G��x�8E>s^��k��F��~Z�9��uN� �h7g��o%����K�����(h$Ɍ��5�ވlp�Պ��Ϯ5!���U:Zp���χ��l(�����y~� 2���Qp����x�0#5m�1���R�苃>[*�S��ۻ��r4�ж���*ݏ��9�����[űL!@�n[��$����:V�mz�a��C��Վ�±�+�-
�d/�R�%�>T��� ��*��~H��]`��G���Ƴ3�Q�+�;;$B��^�M.O����J�d%����@ �����G�=5��12�:�:k*��˲�v�/�ހ��)�~��H �3�7�+�����,\h�����7�4�	����D:���@�d���v��&�Q!��ф6�D�h4�ַ?o<�t*��@�ov�2�z�[��Jȵ�s	�&5.ŀr�Nw�$�\�����*V��wR29�|��<�G�G����^�H�1�c��:g�<�d��*�.��^�=u�{�f�]�T��0f*�	9�9�<ٰ�S͙�^���)�Z�*k�(�����˵h�%����i��PB�C;����t&O��z��q�)�L����0�K��bg��R���S��7��!>,���Kw�.M6A��7�j%R���r��z�`P�6�b��#m��q�%�����W]!�z�(J�Z��L��ؿ���;-#�����W��nv�EpM�-&��x��'��=�
�8���F������c>�R+��J���9/���ca�H�E>@���KG
�˼'V� ���\�z�������η�c�Z�6�]1�d{����D�X�<�>o��*^[%���,��-�k�����_q'�X�	��F}��>��SJ�\Em+��6$9}����AΖƚیb��fȋб�_)S���tLYȾfu�*{7���=�]l�B���^ ������C�4�KQ:l�Y��e�A��CF��c!�'��M�LM�*�ͳ��=ba �S7�{Yצ}�AF+zÚ?�2��9�1�^wC�=d�k���:�K�L~ >�|����K�mpF�v
���Ҁ���M�'���Y��`�����m�Ui�ie�@�<:��x��RN���b��qҫI��]B�J�թ���	S��к�z@�7efW����ț����݀]�t0E���Rl�䆷��1��;j�6��'�z��7N&�p|����{�Da�t��]�Ma�Z�h�1@779ܿ�N�+�k�mZ�3&|���t8o�*��Y`��݈A*�)�Ѡ��v[�v���q_�R��I=%��+�K$���6&�A���K���8Z%�Q�bd2��U���/=�g�$�#mߥ,�?�����E��a���?s�ݨe�O�z�g���*Ìi@�)mn�hc_:]�z�q�4�,�O%�#�2�:��G�'ס����DQz�T���T��v���r6����n���l:o���Zx�����P2
Uy�ߌK�a�a���㾓u�ܽ �
�����N)�k*7ƄJ�!�%���m�J�Ot��'�TNiz�!�-���٠��L��X�v�
���4<��Ae4,�ߵB�~,R�S��Vju�.p�{��A�0�a`�V#�k30?���F�/8xV�(��4py����K]�GvC&8p0ا��tj�P�Q8*	y�iܷ�#�C	��!K�Jz�'�F�Z�4kh���'m��Ζ��{���|Q�X�d��>�=.��Ȋ� 1&�X�C��e<Ly�0�c�'�3��/��g�D/�\q/ᕹX}�N�
�,�����u�R��b��x]_����5Z�g�s����x����i��H�I�S{LD�OFI�ȼt��o�И<:���%�4nW�(�!���eȱ���X��ݶ�2))�Y���'�ߗ�g~�;$g}-�ئ�̯T��0m^"p���}�`�r��T{��j9�Y�c��������N6b|+@�wDem�j�?D$��c�2�R4I���QajC5-�c���QP�oj�J�� ����6��s м����D�y����h���;�r�Ag�Z��(nX�;�8�
��4�t�j8�V;�0?W2nڳi�)�Ev���`)��M<���;�z��tR,��"���@�U�_�W���1��q���>��)��va��c��GN+�P�	_UvS���i�#$qEpK�H��|�<Zɠ���f�T$ER^���6̮D}���b��f�I��o|X�a"�0�T��7�_ܨ1AM���#�$�+�.�uUwӜ]�]�Lx$/��1r�qs�"eK6���H��4�3?7��=����PB�8A�Ȭƛ4i�^��K�b���ʤ����V�d0F67y��|�Ŭ\L�JKcZA�.���DQ'1 �\X.��	ڊԁ���ͣ/�� j�Js��{�����0߸&�� ����S�s*��q[�r�S�D�Y9O.�����g�M�`�GŲ%���@��,���mN�;�������V}D>�Q�d�i5@ĪbК�t�u��}S�I�1\� RD:�V��#^`o���OB���^<<L��?.=�tԱ�-5#E���KF������Hr^���sn���z���>*�����Jn/J֝S��8�V�1!g� ��ȑK�ƫ�o��4���X���)�~(�Y߱��/��J�H����W�=R���݂w��LH{r٫���?J�W�ufc�x��- )�"D��4��i��o�"ܮ�����+sd!��7�-��D+�#�P�����d��٩5s��{Đr� �ې �ԋF�P8�1r��Q�H]d�YH�7BW����>O�ә�\v&5���'�+p��X��D�Tg�mG<g�7�6Ņ�W��{��?�bK�����W1���E���xr��{ugOD@>ܽ<-�X�1�%�9����x��Nl��X�Ր�g��{�X���ـ��̻q��� y��4�b�|�%�O`:�I'��:6�9���D��z���ڈ����4T�|b�۱��Y��RGv�#�Ms�A��X�Xf�]��:0@h�P}���[8'��=����=���[���� 3�=�"B��M`�.XX4(b�lD#H�o�~���8:�U��-����cgӛ�&��� xI������{ua���e��G�x�RaM4�Չ���v�MM�ED�'P�iC������kE�dέ��N�3>���:���.���4���'�b_d�h�
zʄ�x�n��5 E�&E��~�"�1د�+�&�3��
4��@Ku)��`����������U�����*����צ�	c���w!6� � L�m&����h�]���$z���H�I݊��_�a��=�����|�^.G���~����#��2�:�vS�4�۲�*�	(~',�E^fpuaʝ�@���w����[I�6�T�N���0��n(Lb��<�5���(��dW~1��a#o>���A����7�ؖ��[P�x����.��=]J���lc��<,����B�-�Ӫ7���hK�Gw8����g�+���՝ĵ�{�;\����z�5�� �׸v6�/��.�TEeO�u���v�fW���0̵V�s���]��K��p5����܋�  �TC������!Q�È�L�X�o��#D���K�\�`0�h��ҳ�`��Q!1��8\+�i?�x-�se�:�ˑ�W6�ؒ���x���'����ʼ0���&���>�bb���"�_Zo��O.���P��Ԝ�ߥzY��^�gn��%OιhZP�`�|^%�;�zZo�ם�..,�c�<���Y��!L�fS# D�C>w�Zs�r
�rؑh��z/��@�f�1�m�uji�]J*�7���	~�~�ῤ+)�[C.��^/5Ae:�In�+7!�c:	��C.g��G�$ܮ�xXޒ�t�4x� ߮@ۭWx���;���9n�vo}�J%pkPtߗXg;����j�{���H�RNp=���o�1�Y�%mF�/��.�0�XP����t{y�� �.�	�
W��s=�}?L4YN�1��	,wY�Pu���.��j6�Ӿw�~�sYw.���2۹����dw��}bz���LkA��%W�euz�����0��Dle��~�>HF�,���&�榨JmJ8N�ɋPQ��.ó0�c�-�hj����,���)4�h�^R�Nz��wǁmJm�u�Ȃ�t�ڇ�ޔ��ymP*��-���;ꢁ2-�\�JL�r>�Q䧭�4_k�����y�v�m��!0f��d�(�㫱t���N��V���/�X�`Ü����V-�$�tyG�׋�B?�����ڪ�����F$[�1!��f��}��z�/.�R�8QYۨw4�r����Bq�N�ҍ�.�P��L`uOU/�t������ddPH�D�`���� K�M�@���Fۍ�,�IT�%��H1�5d���%��h����� �!�&\
�Z�a�n�+�
�j�ICi%p�}q�kE�cj�4���ڙryR�z{Y48����!�9K���<���DP?��x���c[e�d�(`�щ/��<�%L�ף}�X*(����b�Q�	������Z����㵁	9�������X��c��� ����L����֔_��?�$�w�I��l����s�W ˌ�"�=��JԷ[A�d��;�\eݪ]n�	o/���f���K_�J���=0��)q���t
����|�T�ka���~#���}�׶O1�&9�J��k����%�w�I�+VeU	�`N6�U�)Ra�=���	l�Lz\��5��e AZ
=} ֏���'�n�UXo��y�2Y1� V\���ns��[��.�*����0q�V���0��ͼ=4p�a=U���>�&]�E�l��4��p�A�T^*_Y綹']�!�/t	���&��}jH��He��(�S��[nh��h�
�y�N��lbyS׶=��Li�@z#bASV��yLzt��V���v�y�|13�Jf���{ݍ����z���Ӏ���U�W8jа^�����-[����L��[^t?JXbO�2���ƵˋI�$'?�ӏ��esq�)Ob:/��(�������
 G�X��IA܄��k�q�;A�-ZMf�<O͖a�tP��D����D��	��=f���x#Ԕ�(�-;�-�����剚�O~n��(����R��H��QI�sGf��ʽ��pag9G�a"/}:U���
k�W�|�Bq�kC�	6��&@-�O��+1��T��/���ÿ�Ѩ�m�#����7��W�y�\m�����ҰǏ�^)��R^�/���Lvn��YN
-w��Ƨ�����wt����`��=�_���x�5�\�}������`������2��Xw6QwE>�|��Y۹B.�_��.�6/=j�/�����{s�6�=��xC�C+�.�� �1�h^C���t���v��Q���1?�o�/|L$�BO
��[~��ޤ�n�����4��/�m�AzZ��>$Qs!]|�\��%d�,i�>�V$�Z��G�3����E�B���4"~�nѺ�kLTE�}���A�).��9EM�}���y�p��/�^��6xN\����&����䡧�uh��-��S
��x��`�t��Y�L�Ѕ�?~M_��n޲lp�I_X��7�p�X��w��s}Yp���}{l��˳5a�Q��0�H��̍�O �B�Rhl���[w?�_��4���O�3ȏ����urRh�;?ng��p�:L�b��o!E�Q^�r�J����G֚��|W����$����hh�f|�N��X�e�7(i��<L�"і ��s�����?��jz�Uh�/�����c����Dp�G\dg���/�]"$\��%
�S�$oTe��{0=5���$9���Wo;���k���B ����g��"V�XJyO.�?c�����H��m�B8h`�9F�9���VG*�|M����S��@>]��p7O�a�3�S��@���/�)	*�./�e@O�����p������XlxVHYEB    a278    15e09	�=~�Eb:*����	B	�RNv��c)>lwb���}�(���E��fy���&��xz���'�A�~��r,���4��q�sn,θX/�ٙzHlL[�t8"���\�r�p�� ���6d�?�tk@��E#��Q���[d�{	��p�%��[|Z�mӴ����b�g9Q/�Ux���4ʆs�唀\�I���S-��
ڼ��k����k�Ǜy�@�k���y����Q����Pڨ2�<96ux{��ʽM������S�b����$8��q�ys!`�9�1==��*ͬ<𸈶��f�L8�C [�,�2�Q��!�w$�Fq�}��(�����v�J��|ݥ���`o�&��tR�u-Z#��u7.S�� x�W�M��k��I ����eJ��B;���j���)���vtnRv	��IE���n����΁�;HAu�(,bJ���nO����eBui��
&�+�W)��5r�K2T�@��g�����ES}�E�:��o5��Seq��Og�7����k���߆�v�d����f��x�>�:^b������������S�U�Q�&���9��vFE2M����Mk`�+5h�h?d���Z��A~���e��MŦ����F����2n���E�Bi��^/��}�T&���*�c�ǿ�q~e�1&�DL� ��j���S�'J�{/�̧��l+������Jb�c����]��7�xTκq������� �lye���Ə�(gm�Br�)|�H�D�"h"���-���j�zǊP�6���j������$��!j������+E�ޓ7��yUj���J&:�z`�w�+//L��%{�&ِ7S�z��k���,B|m�R)�������S� ����쬹1Sߒx�V��u��6�f���W��v��f9{c�)@@E�q���H=��.��np�� �O_����� �뢓�׺9�&S�S(����+�H�0���n�i����Q�<��q�G2J� �V;2r=��O�"-kz��`z*�I���������4�|��b���UӖ���g�4^gĕ2G�q���>;�ude�5<Θ?U��Ӻ��J��R�r����;F�x����+�d�c.�Q��r����A�D��79�ۨN�XqELڳ�K� �G��Z=DnC��� ��Uݶׁ�����5���r�YӖ���~��܌ѾT�Ɨ=��LN���=��s?F��aPi��[v��OsZj�X��S�P�GȖ		)((Wvؔ�=^�V�.Q1ʡ�#�T���[E�B9j�q�,}��e��u�6�Me�`C�z�,^^�LE��
���zt%����fe*�1ƌ��C�r6��)�U�D�Z5P��?��\/ �����PX��c+_g�}��B�%{�7���Q��%P�5R�|YP|m�,٘t�Fx�ӕ��|2�U��u��|���$�vف���{<�8|Tb���v����E} �n��#&�v�]=��+p�0U����<~'<��*�u�-J�:�wMR��g�Q`xR� Y% Q�n��b���+;�k K�6n��fj�T�E���(�mSB͇�X�o�w_�����/l]�Dc����,Z���;�~F��UvO�5�E� �p�'H�5��K��D�<N(?�+�Pއ�q@�P�}X���^�pݫ-�����%�>?���-ʐ�$��|�7�%Ρ��K	�%��= �0C�>.���NI�Iu;���~h�p5��<P{�kt�-���7H�2��w�Q�����P����Z��3s��
�2��vy�Ӷe̝�J�6�p$�1�����h��*�5��b��nQ���7_�	��������݄8� &�|/Ƞ��
� /����
$�J�'�"�	��*�Uf5K~�QƔ���r����5 ҕ�����#�`�Nڷ�)	������	2L��z�G²�J�P�A��^���,4�"�|��w("�C,Ik���FBA�������~�dQ�!	���Q)P�8t�����`x��Ex�8���>��I����#^��@
�@�2��~w�|IА2��q>e(�����3����(�{,��Wj״�Ma7VG lSA����2��q/�Y��}���L��2x���^���(qi�������n9���h���h$;��P-S�dV�:�#���X���-𢧖�@��2H\f�Hʃ�bj��J�Dn�1�[{j_�</Pi1��1��j0���JOYHb�rQ��I�r��61SwK��c祜��0��z��k�����K����,B��%�O�����n�l�;��'��ܠR�DĆ����>E��40��B��78���IW���UE��	���O��Pm��w��ai�j�z�B�w&��}�� �e.$�bUvb|����C�u��1�ؙ��1.Q6��e����V�%��s��
?M�J�%6�_�����W�o�ђn�&�	u�������h��`�;����StE�x`�΄s�c3�c"�	e˴.�LJ���O�N��@Z������<���&I�� !��!zm��� ^4��y��÷���,�����c*�gv�U/�)���� &iG,Z����^]/J�˟H��d̞A�صG͐�$�HZ8ƅo��p@�R6U2\�_�B9MLa����D��T�gdw,�ב���۰�Z�\,������{c6؄��X�LK� �e|�
��b���C؇+�ܢԸ�-�h�
B&蝽��C��bP�9�PKRa�������ؽ�(��M"�m�D�k�[� 0���$i$1�k�~��������f�VI���A��E���gׄ8ɘ[�Z�A-l�P�hoJ_j/~�S�	���!Qq�Č��>�)��m>!�ُ�߸ϨD?��D���	g���V��*�`N���2����.�L�M��UXF�n��<^�uF��������ۤ�7y�� wQ��Q�A��
�|3�F�G�]X2��L���R`�w�M{P�_�ؿ=��P'���.8{������r��[�?9���no(�qG��� �b<�QwR*>r��Y�#�\���$e�&c�w�
S��d@Aߨ<ō[�#gv�s4I�R�f����.��d����2��8����#�hx(ި��8I��s��n�&�R�?�j��)jiawм^uߍ/~P�y���P�n������v�C:J� �0�6UjpRƕ2���DPn�����P��&wEH
��$���F���⪲���>!���������L�M�����BLhӅ����#�q��ٴ�Ů�����N�!p��Hނ�^�p!�g��<�E�V��_@�P����9^��}	9��n���:�<_���$���3[�c�q��ږ����ÕBJ��d���`W%=Ԝ��W��I��daP��ܝR��_-'"��,�4�3ŝ+�ެ�lx�h�i�z��Ͱ��t)�-��{w��wy�;co���X��6{��!c�R����w�h42l�r�� lt���Q���-/QS0V�1��iӶʟ���"_+�L�H��<�;��sHc@�/p�[�뉬
�6\G��瞑`؄�R|aո@}*�q���\8��C�K����]�8�C��CtހYP�fS�t(����=�$�@F�,��g �<��7��de���ݸ"��+S��jbz�׋�v��gbB_u9�tR���{	#�&���h�7�\��S"\����I��F���&�3?�F�
�ac)֯��}�m���N%WR55'����$����od��1�J�l�	��ɾ0K}0��������n/��v��>�C�6�z�l4^�Z�T�kɾb�L��N6���:��qG �Fw��`3z����0]&z;�)-�j��RY��G�&H�cK����	<*�k���3���.��%�ɽ&��0歗j�Sa0�J&H��Ih���Zk˨t>W���jYp/L"�ڌ�_�PB���*3Y5/�2�!߻�q��D�A& Dj����XfK���'������0�p���8�����$*�Ώ�e���G��U1O_�:6�B�|r����dBt����}�BV���K���j��B:֋��bdݽI6�'�
�N�����)�r���Q%'dѵ�p����K]��O��$��A��P�Ei�0v#e�b����׻�Cs ����,�y���M��al�+���^��%V�!�Tȡs񈨒�nߴFx�O���]?@J�$]���}9o�}���~U�K'z�ue+_	�a�v��&"yZ�m�AO�M��j<�i������X
�DOILb���<[���������we��c�� ��1\	-͌��D��V�Y� �渿��o,f5�ǩW�f;{��Ya>������?�.���Rro��e��}�}��aG�[��(jH,�����\��+H +�7l�0�q���q�g�;h@P���(�&6��1��Y����b��'����:�J��h
_8�ɱߐ&[��0��v4VV�p���M=J"��`��ߍ�7�d�S��k����jL�<������w�!:*���|̢�S�*0�: &�B��_5A�9a�)ըLZNU��g[�&[���|�:�l��R0A��S���*�2�$���ٍ�/r�A�_�X�N��#wrx0]�_��Z�>}"��z�Pl�$d��������G��(͸n�3�D�����O�u�$JCd����D�	NGl�l��[�����b3=?��s���N�uj�F�H]��'V!m�T ��ss��6W���g-����vo�C�yכ��"��E�=V#�y쀦��� �r�s�TaƁ*g�+��<��Wxw����_���pɥr���u���Bbwj7lZ�� ��C2���m+�Uw�A�'	+Σ��%��Ku����24k^�c�i�Ļ����94��\��>�O�l O�
xd�<��S��S��#v�m�Ԋ��0�L�=�W���E��1qZ^/ւH3\���Ԩw�Y�HW9�58�.c����_��ʔP;��Ԯt:��n0��(������_��p�p@l_��G��2m�i��3���9H��QCF4���.�)t��L	�u���ք#�Z�����7�?��W�	�l�[������0�������!�V��\�?��gA��Pp3_o���Ӊ��Y�nV��eQ����(.��YiaO)	)L5�ɂ� MU�������e]7����s{<K,1��:���m]�j�����:*Cd�
�C�*:�BS��7�� ���vhN�%�����9AWZ/���RpA2��y�p�K�����GMZ\����<p�sb�T*d]Z�d\�����m�D���p��� \x�p)�[˔04y>
����C ;~ue���_�	$&yz�&���m)�� �%��I$�3����% � p��+�,I0F�}�E�ԃ&�:Z��f�����Q�0��մ���
�7,O��ڽ��C�w���2���6�����