XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��qh���0�h�'�J )�I�k����UK��u�Jb$*02���Z��Q�0Y|K�LuQ �*g���P��� ����*�[=
�bS�t٩!�2oE�#�h�א�����n���΀{�<ʅr�A��vf]� ��)�?���k'Um�Ec)�9m{�r�$�;WN��~��������6��b��2�P!5P��?	�Xi|�0�!�2t�T3@�+�(G7g�u��r�A�^
ŶE|��y;�<쓜�����l�p��Ē�B��n~hZgtq9�ǰ+/�5Ai�hJ˶]�͚�V�P{��+˾ӄC�X'�;W�����v�,��bֱ�2��$h����1H�۫�∨
����Ɣ���R���d`C������J��h䗿�zs�lj �|p�9�P���<m �
8��@w�*\� �X�2�$�^�k�*��:՝�w�=4�n�����Ak���5-�x~�B�#��6�ҋ.��A9�F��GE�@�8���^��U.�aVx/�X�*6��c��fZ�:߹�[H��y�����������"X�*r�A�]��.8h�Mk�tP�>��9�p��Uښ��r* ���e���5Y�ڽ�З��������c} ���_/�0�C/:z��M$��h��~�i���m���"�׸k޿����5^�0ވXV�o�xυA���V��y��Δ�ԇd��Yc}�2���(�|!�$H35��d�P���ҋ���T#u�~����";ɥ�q|�XlxVHYEB    9fc7    1fd0Sd3��#�����~�n��W��^�|~��3���+�T���ڀ/�5�F[�����	�,y�S�'ֵvn]S9���k���-���BJ�-��-L��A��2k��!]����}�>�i�%tE6~�e���хT7B����7o�li-Cm%EFp�������[C,�%cĿ^�u����A���ͪ��0U��c �٧\���p�C	�8��F�:���Z�>�0d��V���K����|���|���dp�V|f�n�E(�<%�vz1%X���P��Rp̟X�V�&����S��;jc ���'�9Iq>I߽���!4�wogфCG���U1ڭ�O�
o~)�V:��r����&6I�B��m[�MY�*2�f�e�Ѷ�8�}|T~ه���	�>�)��h�U2��:�)�����nؘ˛����K��z3�"x/�U��Y��ΣC|�4�*P�;���޹/��*$�	��mf��>��t� h8�yj���tv���5x�!�9$���07�h�X�9}Ji?ڹ���}���;,��h/��I���#��DQ���I�1��yn�h�`i]k���
NM���Dim�@�;�
��� �6�i���g��
|��0+��� R�X�)ጆ|�H��3�y"��L�З�ط���A�	�5��>3A6�*�W��C�K1���xA7��N���ݼU�G2�_�/����E�𮒠xNjy\.\˶$�^q����NƔ���{چ�$�z	6j�~��öC��m�G�t2����L��*��+\�Z�>��܂�ZLf�|���VkT&�2B˔-R�/�6�$a�.k���,e9��ã���Kh��c?��{7��=�%�#�wN粘���^���,� �_��Ki��D�Z>;�O�q�G��{Ɗ��
!�TI��1����)��9u~!�o�F�~/,Ѳ̀?�K���B�4{
Cӫ��g��=�!1�g���[�pP�l3iߞ�W:ra�
1^������p���]�W�zr��'3>�q�:���Q�}�@)�
������>����\�V����@{O'�b�� �'�8��w���On�أ`d�*�AJE}��e+sG�?B�_5��A:���C�����0�!lK��2����t����� s����t��H_�g�u����m���b� ?o�Ad���hY���D>S���q5��W������ 6�L�YX�,%,��<�m�.�E��Ƌ��d�Sѥ���1�'�Q0��\J��t�\��e[B���>�2,�_�'����Ik��u�ڈ/���m��+m��~�NDj�����8�Q�(�Z�iGڹ6r}]�������p����6"A!� ��ba��w{��S�,�#j�e�l�d*�wK0�B�pl�n�����Z8_T����#?96�lnf�v���Bk�,��ۻ���_�ʈ�?�b�&�q*��E�X�D�4��bfRu��L��$��T�aE�|��J`E�3�c
\Td�\5K��H۱irh�Ͼ#�6�d��[����c����=�h��-����\�ホ]Ǚ�:9Yl���!�ט��>	^'6��7Ѭ"H��6���/6(�aN3��8�Q��Y&(++|�9��U &C#p�����7Edȗ�9�xe��]�8�y�SR�TM��8�PO}�'%ߟ�W"W1r����e���|h����&٭���+OF]P;�q���}&�e��UN��>��s4���$��Q��1cc\�|�uɚ+r�����F�h��:�1ְ���>\!���eZ;xШUR�����
i@\�QMl�X��N�
(��w���?��c�ِ�!���,y3�a�d�$)h��τG��V�B��Q��nۄ�N���d�	o�ɱ�ENG`l��oU���Z�L�IHaD��W�;��6��A�5�A�T�\##;�Q)�kRyh3�a"Z��`����>�"�m\��t��WM��lZJ$j-wS��#X���[k-�9�0�٘�������[�y]���=?�K�o�̭�>���"�<�uWv�����5c����-��W?/��Ǘ���=�'��|L��E:4¡y+y��Dг�$bw���M�(�9I6�L� �\�§�ӡ|{O-�fE�-��%!V"���-'i�2�r���F
j�	L0��]y�,62�Zߢ��U��R��y��1�*2&m�C�5�W���%�U�pP�{B����$�j�����<��w�|�65������w���u>�cV��"9q��Z����A9K�F9��e���,�l�F�)���0¡�*����+���0g-�X�8��$Jv����谕�'F���a=M���(��_]�Lmmr��X���2�ſ<��I���xWK�F8qn���K�.�׹�K��!�|)�W\�Ph�j$ŀ|��1�s�������������j(���]�.����m�O�2P}0-�z�$я�;�2 ���0���f-�x7w�#��^9�zYh2k4^m#�;���ZH�G�$@n����]�k����C�T��5.p���s��}&6z��&'C��!_r�����i �/��*F��^En������e5f�}�p��y�!cnQ�؂���ggǁ䳽`��;�e1y��M(�D{��Ȩ|��c/�q���!w��'�Ô��̇O�r��m"U��5sQ�ᥙc��`�$\����$`�]ǩ)Va��?������v+�Q��@����*oƂ�xV�"X��$�Bno"�;r&���XW��XU>%Q?�if��܍��Th?�K�vd(G��g��t�,hG�0��b�ʠMC��MF���b���o�o��ʬCM�'Zd]���Pb_zA;y��	g��>I�C�&C�M~��Q�*���H&�9��ƿ�vU5k�Љ�Q��� YH���h���Ϣh����A��"��D5��K����e:�F�ImF�>&��љ�y�������g�\� 'vj�gvF���n&1�c+4o��ͽr��,��B���fӷ��6��J�bqb�nS�+�P�<ʊe��ҡ��O0 :;5�ɞ0��t���	�*B�{~��D���<C��"o�
$���kE��2�
:u� ®��G�^R*����t���ZP'M>�8��V�v)[ɽ��>)�ˣ= ���y�$g���Y,C73��zۜ����q�4�ƙr��p����e�
�Pް`O9k�xs��皆t�L'�(��L�[������ދX�#$�~�Z�`65������u���/[^QctI���M>0	t�#H��4�4��{�ٌlkI�XaO ������.듃�����SP� �Ei̝L�)1,�4Sy*-6Nх��>�7�����T�[�_���K*�E��"�n��{6�B��6�Ƣi��J���L[o�2��(�V��qa|�Kj�.r��w�b8KL���\p�������h��}�����Wrs���l�k�3�M��T�:gb���~J3x.��)y�T�x�R�W�g�0����=�wg���3aj1�i��R��m��H}��}���'C�؎!�i�@%pNY�4�
�GE(�곫9K=��j���4�Õ��ƶ��������
+P�z�w��6l�K�S3��) �����3��MGG?hQ��˵EvF�ٶ��X��G��ܣ5F��������aپ �k�T�F�0�����e��(k��ρT�j?ga�{&&Dm)G2��z���S�cGC�4����E��Vz�*
��_�����9�S�K�ޕ_eq[��~w�6.�{��=)(���`���~��k1�n�=��/���?���#_5ItkT���t �����U�`%�K^��Y^YB��!�Y�蜚5�J��?k���H =�+���m_����^N��)�_^��$?8�&�Gv8;e�˒浞�x�W�g��)D-\��%�] �]p�Pl�.A<G�W�5���rT�̭n(?�Zs�k���l��Y��_����3�����A�*)�Σ�v$��7L�<ީ�o��p�eK�����\����ѡ�n;�N�5{���qa<��:"X. ��Z(7���[)L�S#��/w�ԇ,�d,�^=�g�@�#����V�����pp=ߛ���U%PBnΡ��{���ۿC�B��f���}�Q�����kS�<(6^S9/��͒ꉦ�G*��س{��1 ��F@hDl+c;���x�t{��&�����DL��uhW��"\�D�Fr��<������;��= b-F�F=��5!^���4&E#r��|�l'8��<{+�p��+�-���}E*���78�+�F���;��'zL'E��_��{��E�����y��4'-p�;�
+�:�U<=�l���	a�֍A0;�̃{Hq��N�b8	|�k�6VrFe�N5r>o3'{պ��DD�8������7H\s�R£�����N����'*���_H���@�3ٺ�Y��Ç̤��ٸ��s[�t��o(����@aJf���S?ssw��>H�b�q��Ԅ�{���l>�����|k��/{V��W"���(Z���Ǔ�S���${���V�Yh($�Ά�4I=�;ʌ��]���F9B�t�q��"c�n��oe�� ���U2(�;{u�Qx�^�DFK�r����Xh���g�	�\>vY}	�p^v�����.q���ap�U �Ɣ�j���C�Bɥ���U}~~O �*Ԓ^��z1���<��׹R�`�=��>k�ϥ�7���H'g�0����!$��~�+�x�C��(����S��D���`��i� ���CP߉�֫��<#��Su����
s�|ջRw��t�(��T����\��N4��&!�����ȉ,�p�\g��A�U��O�x���!��K��6X��,�g��d��;�i���}&d*l�	�פ{5��$�9"�֐�>l��֭��0��US���O�@Q"��/���9�+�V���)Q�&t�x!]�5��Rn8�\P@���p�W�Y򟾲�_8nM�E��*���D��"�e� ��K`:D9��4e�*>��ep�M?FNȱy:E=��
Rs�!�B�f���e�T0�^�P��%�s���3c�T�!n	4�}�Ɉ���j� �����ؙ}����)x�h+����]����g:�=b�u���fS�<�HJ2�>?�l3����`���f()�M��	x~9��`/Zst�� K,��*�%��B~u�a	GqR1����ZB�q�4����_�#��
�HǤ������{Ҡ�[�|XO�6�}���{&˽2^�+��t�� ��l�-��R��pXk���4�_�;~�/}q��ʳ�U��q�ͧ�Y�N�Pm���<*�V �Gf�ƍ�ÖI�8����B�[8O���"L���C�I�g�NXMEjh�#x�n��"x�X����ܞ�(�d����tl㈔z�Fc����{�VVG���'�\M���#]Tlr��s
��^+)��\5B��|�q?ST:���F�k�L&��pN���kgT�a�`C}�����[P��m�.�V3�I��L#��~!�-a��SǏ��W��ո��	���a���5�6�tL�f���5S*�T}Q��]�2O�S"���5�t$��6	��,��o�o#��e�54�[�Qc����<G�k�Oַ%��B;�y�l'�ZT�~���|��y�ִ���l�^��y�ѥ� �Y��CDdN�����ۆ^���7�󪚉�$(n7���3C`O�I��F�W4w��(����	��#���k2��؈�[("���A����O:{�����Z5�֙��Ota����C����It/&��ޑO&Nb�p�;���}��ڈ��\-TI����BYa�y���Z�H����v��Eő}*u�A��X淠��$�q��*2i�[�E%�� �>�zfB]I��K�q��]rd1����������0&;� �50�0��B��y��{��5��t��@����,���Ρe�����8���$ʔ�{^U)K�C�m���c��>�dj��a���i�a�COs[��z�Q�6zB�g�j>�J��q������j�^����[�����C_�(\"�E������'��f�\
�zϹ6�������������JX�0J���9Yus�
|0ۙ�D~�w#�ޒ:_�3�U��d�f���r���+�w�xM�>�>�.��xS�qQ������h�#�'I������Q�֑�` �yrH�����r��<�ь��g���.&a~0a"���qY��A��Rv�[�~
��-��U�3���H,����ʱ1�qQ�m5�\õk�.-����A��%����<��e��c#Ku�.��S��
�=_Y�3L�d��:�,�4�s���(�+� ��5���)D��5�&-V���Q����)M�{��+SV|J��P�reI2�pGI�����8�*���N�r9ǫ���Ap��ҹo�/��&"��OvX��o��g��?���٘�ӫ�2¡��a�@�:՚����#exY��U�K+�ƻ5jò����V�̀�}��9�F�K�-L��U� �HUC��`��y_���Xf�E'Vu�J����L��=	���hY�6�9˙�Z�j���}C}���[��;�S	͑c^,_���_Ι+6�+�=Ί��h���b�;v�6Q �n���#�����fB�Y�#d�k�q�U�d10蓅���E4��u/�s���dnLT(�(�*�Ԯ��r���H��V��k 4�h�:����y]&՞�v�⯔�I0��Eq�ƫ`�I3�wc n���@�C�(<{�L���箖���3�Ҭ�N� %]����@ZFO�c�͜�&�4@!�7���>��GO��}�� �	����'���D ��� ��\�m���|��m�g6'�-zϮQ+�o[�u{.g�m~�_Q7@٨��vh���R�5 ٔI��b��_	_L@�=I�D%P]��CR��YN)傛��-T����Mĵ�g�71<?�Ʉ6�pA�=�}��@�4䞽�"�N��&(����!�V�$]�VW׶7S)�˘�,M�����$>\ӏ�U��J���s�E!��P퓸`���cQ+y4�8�\�����͚6l���m����}��D*�C*�GjM;d��96�3X-����f�Saj��_��,. �YV#�����m�O ��3�=O����k ���ua�lX���n�۩0!�:[]�/�����:F��\�r�-e2��k/�b��6���x�^ �0%��T�ބ�#ݧ��djV<�T��x��Q�ba�JAg a#ۥ�w�$�ޮ�قp���y.W��5�_͌��/Vkàc�T���gA��pC��0�Qx1h�kv?�4n�دO=Q0��mm�#� �ָ%ʻ�a�4��1jGW��}���J�Vq�������_R�8Y�P��ެ80��J{ ���
I�3��c,��r���w
h���/6(���e:�?L���:+9�Mg૥������;��S����I��
LSM�u/������Յa�*��������M��|.��$G�52��6/��>� � �Q�{���7;r.fr�ຟ"��.ٛ-(3�-E�'u<��y���6�_����ڲ��#G-=���@�����f��z��e�<���]�_�wB�r�4��,��.�0��w��Y�Z ��ז�J�-�|d:��~����q��U!�H��Ǥ۩�.�UF��o��~v��S��
N���c��%�:JE�<*Gz�qE�"�~�o��Y|��^'� W�&l̨���pt��m
H�B��)!�5VhQHT�ɽ�5�39:&�u�U�ںL��fxUj��{E���a�V�]qޏǏÅ_��E�]�,5�����n�?3�8��/$�$괣p=E�V���j\�5�S���^��w�ť	0P��]��[�"�����bK��Y��+�A+����A�Ă��S���
�C�й'E��6��d���c�&�