XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q֒���xW����.�q햪�:�JS�%*�;�8�������K�B?�躉`�1�����y�	�1e����ǂ ��^�	@?���&9��񧣃�KO��^ ���0:b��ڄ�v8Fs,����dH)œ[���J�g&:��HhPa�T�?mU7LL�_PǣVE���Ց��2���|
<�A�ǒ�� �de�f�T	��pQ��v����T�{x������]p�W]EcX9qΪ��Y7�q�ӻb#�u�U��ݞ'�^�~����v��\z���S�L��^R��j]�|�-R�ȻW3j'DQ�H�L�Z3�L��[~z�r�6Q����j�]��������v{�E�ȃ�=�%�I�YۈT	�Q�o��E�?+;�"(ҟv�V�I���C�m�������X����DN�P������=Y�	w�@74X�TO�>@��g}����\mv����:�.C��潆�M4F1;��w&��?N5x��N���3�off�������%�\{r�Rp�%ۖ%�W�6޸�4s��8�T���6F��>A�a:+�MW�ڿb-�������2t@��8E����U�Xod�A=�ʳ�[�|2��Wl��f���8�ZWe������9{�~u0����1��Q�f)�eŸk��a���Zŉ�!F��[k:�f�D\�����%DB����l��}�'�ζ`e�v��� �K7�h	;E��Y-c��c?����u�[-k}��;�d�s+27fxq�&���5j���+�XlxVHYEB    6315    1790�+��x�t=_�+t\�bKYL	4����o�H�т���*��3��G��T7�f0"�V���	!!�����?��	IxJMb̏��d�k�c�}�^j��u��ۖ�I�:�;��p|i)zU�Kw,t��]�#2�|�m|������f�шx}��w�hf��z��l�I��!?W0�*xvn�V/����2�*������y�S�#��M:ϩ}�����
��L�Z�`Z�I+��I%�i�{F�Rr����-SVz��$PXO�~ڮ����O���D.���������j����q�ip����7pL���ŋK��CV����hh� ��C�#��ڐ�)�:�?�֫�<ƽ���y�^��_��\	�e"D��Cby�E�-�������P��exT9�M�����ڦ&ބ	{��Y��*�A���H����'�_k�`��Z����Ȍ�q�'ž�{�5| ��1X$R p١����=!��%a��Px�;v�
Q���i��ͷ�	�}ѷ=R�k�#z��GR���]o��(-�3l���I��e�@��1�'oU�+v�0���c�/�h"%#]׍+���|Zq�I��eT��+��L�� ����HJBϜֻ����BD<�G� J�S�ܢ�*ե���r�d-:s-�3���9W����5�i;awbk�6}�o`�"Kr?�E���7�Y񕘺Հ0֣̐��v��ʩ���x�pDۘ�^�;7�̴p!��%�wj�t)��v�@{�ӡԪ�sab��T�*����%J�rx�i�D;5���To�bMl��|TC�2tzñ�w#�Nɀ<�������]f&H�l�3@N��Ĥt,�D�pɌ򛉪���[*oY�}�b%jY(���6��_xyW�W�t=��1��*���UM:�y,���BC��k݂��y8���ʄ��(�j�49���o\7�P�{(�5k�S�~�rLc��^�(��h>^�X���CLnЭ@H�����*6d�����a�^;��q?��Lk� r�����~n�t�=�*]�EQ�Oo��g	��|��+���b�b�mw
�(�rǂ��&��qO�G��;X�~�L�o������$��U¬J0��t�	'���L�ʵ��ܜq���Y�n&�w�V�b4��X���:e���ۢ�Td�A�c>��\KT��&0�W^�cc,���~��1�����݁:�U:2q���(����6�}5����<��st{E��Q��������)�t@�a��#E��gm�Y�ˎ�e���H�4g�sr!<|�ɴ��X���;pb�ڹqQ�9]�D�96�b�VI�����Ȝ=\DJ��Mub��<QDdFv_�%�����3��[�l��*��p�^��Տ�l���#�Au�"���%�*���*07t`������v<�n��0�hҁ�C�E'���K����֫��z�`��:���k,�l�`�����+0�;�m<=b��q��B�<�s�[?�K.2kv;��/�	v����!6����jh>��9��)�����������a���F6u��a/������I�1PX�	�W0���4j�o%�'�4.��T�f)=�59*$�Ve	���qrh,-/9#���zg���p����	}^�	N����TM��Y�' �ԧ��ħ�F�e]�����Ӊ �� PB�xr����KLq��{�6�K����Qz�0��� ˶��2�O`Q�L�ߞ��8���;։6����
�����MUh���c��Z�>����6�X ��#�gh���p���>O%���p
�<ā��':�w���6f�X�I��8��?O����w�+i���������\���]�n��o�#C*��^V����z��S������y�y1;?[5E�]��u��ޕ	�<P�}f|�C�'j��5��b�����!��(��Z����ĞyYe�פ���c�H�h�&��z&���6ۯ��"��;t��b�V�x{y#��o4q�Fj��P&r�9T���c��:@�F�x'�,�(4��x
:�P3#�O���I������G�kۧ��C�#E��ܸȆnr���A/8��B�~	8��� ̃��?���A���v(y�l֝����e�^W�7���X�/2�҄�0����|��Z ����ȶ�� h+��M������i�~�H-��c��4��J�+q}$�!@�I�J�IИb{'�c�U��\���s�p�?��s����:�-s� ��Xd2}r_��n�t����~�v��.���cv���DB�eVq�ʻEs�\����_��˵Z�RIY��.������0��w�O��}�B���l�}uy�L)t�w�6�Ss�!���㻧1���X ��z��t���x��TF��}B��R>'n!�__�ݦQ��q�	d�^-�P�>�g�;�PX>�s����թ�|GL/����A�t*����F�I0��H���[�k�e^�9�������}l����l�EY�rԩ����*�T�R�2�E����y���_W�������rYT��/pYG�P�,������(N��ɮ��}{pl?u��Jߴ���R,LF?5�+=�6��\g��S�2K�y���g��+حL�f2� §����=�u�g�^����>�4�?I��Za��
�Y�Lޚ<8ͨ(��7	�1S�u�[*�_6��h�ńKl���
$��U�ny�FОv������ݜ�{�����M�����x1W��wg�b�2ԅb���-�n=Cy��2>)s���:(�%FN���D�ҡ�edef���{;�()/D���hz����g��3��a��m��]U�����,w�Q�ڇe��$eH�Ya��,�pLm#Iܾ���\�BIH�����}U�+ ����-�I$�=��5+@�=,](F�]p�)��t�����K���З�tM$�uy"�:jB���\ &���D���w��RD�H�V�;뗳B� l�גS���Z~�:O����SӨ�M� ��V֨��⡴&/}���X+�&b�Ŗ��A�8�i����5n��q�aM�1�>ۜ^M�R��lN��=��@�����?�a?����	ʗs&���c���E3m��N|4�zw�(�	08t�;.Eʁ� �n�����yN����@�d����B�?�9j�8�3�������,���Id`'�>����36�{8e<D�Q#90F��s����В&��(i"��%`�r1�M&�ފ��N�*� \�ԕ�<f�|JO�39<S!7�/�U���Q~-#��xdڠ����s��Ϙ��U�t���=	�i1�Ɗ�Y���>m��(�� ��ECl�Zm ��	T�������#��Nh�����%�[>�n�`��8�֕٨ /�g�̹���n,悄��o/J�z�i�ǐ��1�3,�8�� ��h`1+����!_�M�� �Ǝ�E�uu�dk��D�� 0�G`�.�����TqO��:�0ri^� ��kꓮS>4�BY1�q{�a3�/v/�3B�j��N<�xۖ�&�bc���@�x�^�G�r^NVj�V0���<]~[��t��PԨ�[4��" d�6����B�A8�9Kތg﹍#rR^����� �MP�C��
w�������!�㤃� ��x?l������� P���!�#�j��>|�x�H�����?�_i���|�ކ;*�R�U���^�e��������b�xL8�K?�r��?@F7�`%�2
��w�}�&p�q%	�qK[�fΫ���V�N�/&)ھ5p��ۮ/0C�|�v�W���E���i"�5{]�h��ؠac+����~s�#�YV�Ѷpo���g��!�G�1廉�����sTW�T��o���ʠ���&yT@�Wz:�/L��S+�ߑ�?���Ƶ��At^����Ͷ�#���Qs��s>��q�a* ����tz�V|�2�*�zcBܤ�R0&:x��tDak@��[���Bmu0��� @�i���>[kNM�^-ܙթ5����+)"p���R�m��.,w*��B{+G���,��-~�����5N������)7�P��bi�c����-v)�F��5@K�F�g 3�k2����e�l��|�����%j�J�0%i$�ٔ��X�F���h��+av�8��i�v{P"��Z��	�T ��ܜ��8�o6FJE�����=��3$�A�b�YNs*=�{���p7>�!c�P0��1�%M z�H]��:���X�������^:�2�|�����`�(��k��iD��dȃr]7/�Y�'V`���=������C��P�P�
��zt틅��j�R #ϡ���:�c��.�N%ksG��i���S=,�W�;���* Q�MC�
.ǹ��,^���4��g��[5�P6��N�Mٟ����q�u��s�
&�?���n�f��DB�s@�������j���3�JF��̛��	A�|������я �:��f���n�n�;5�����E�Y=8��&9	�ɑ�.?x��H�Gl����k]*��+�jt���Rzq�AD7z�_�^8��u}�j~�>�����}�@��z��;f�œ��W����k�<:q��l���#�3-@��\-����)����x��<h]��.u��� s�[d�S5�d�tk����$�mų�v���`�����$V�(���8^H+�l��V��
 i�d�%�녺~�ax֒��D�����_P�,�	��Ė$��m� v�*_�j�B��g{�P�'I��v�i��n����(�RG�K�?�J˖	�'�N\�W`�L��Ae�ro�-\	֍퍁��U��Lnyeͥ�g��n܅p��ϯ���$�,�
q� �S���R̪��%�X�����+9S�}:p�x\�_���e��B��d�<��\�,vgi�+���f<g������9�g{�7�Zu��X5�ጎ$�0j�^�3��܆���k�f�J���	��):~��\��'��t����{�xON��@6w�c���
��F���'�C�)��Hb�[q��x�C�b��K�D>�?>w�G����{i|����L+��rkZ�_sT�	B��?�U���@�XUD>v�c�qKUIO�i�����n?�02K�{U���蕰��@����X�ː�g��hv�+��� �x�ܜnOC�[jVp�-_<�_�)��U��{�V�"�	�re��8�}bR�L���6�$ܥy�+{�ɯ<��M3�=��ν��on���}k*���]J(�%洝o���Br���B@6��d����#�(�)��MO�֢֡���$�Z�(�ېKX���^s�����t�]�SX��� ;�n����nj�W��y�HSF��KL0F83T�xؼ�{�9z����� ��h��Ld�g�;|�
C�������\F��G >J�!֥i^-�}��Y+|��O~�e�n9��q;oi�$��k�?T��I)B���&P��bF����X��/KyQĞY�֙��ډ�l�v�wT�`{��`��Xũګm/��~�;�� ͊fP�"�6&�4����Cd���m"x��Κ�10�ck[u��f�����;�Oo���L�K���B�ب>f��)'I��Y�.d���B�ccK�Y�%���γ��a6f�*`/u�gozH1���ϗ_g<���#B�-�X��:P������2��E�j�I	�F&�:eK��*����X9���u�ge�`�gk�{bL��A�@��T~^&-)g�2ϴ��`tC 1,���ri�:��pI�L~��Т��jb��f������n���,AFm�O֛<�;`��T���f�