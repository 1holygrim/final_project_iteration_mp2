XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q�A��F�!�:��ڎ�u�5(8�4���TL<&�L����o�@�3���_쯜��6�)�o�gW��}/>Y�B��a%H��WX�eɧW鰁��N_�O7lJ��n���ʂ��	rN#t|��Q�	-���l�UD��S��`_dL��_�<�����;�b�csZJ�Ц>>甖�uE?�Ǘn��?�A��6����8�7���)����
v��0�#�h>$?;?`�����ő_���?�迂��ܟ�--��/\Mؐf&ɗ�"����J���\>ol��=[�"k���l'A�GO��F���dͽ��ά�XE�&�dȥ�	�v�<��Am-(��7Z����S��z�6OA��;�����p��wȟ���<��� FKG��YgS�~��\	��Y�>��G��O��Y�TT����}\���2�4��sq\O�#���پ�����;	"W>�>��J9�ޜ#䉺T��+�UPR:[z���6ez�����Ο�ѩ��46�b���$�GG�e�7�i�����J3΋/�%dg_���5J�ME���BO��m�態�z�3��RR�0i�>�l,��b�n]��»�q<[H�E���x9�1�0��X�U�Y�b����lE�:)��ʓ��1�b�	.PW�W���P��X����� ��
��r�Vң}���3�jobƑ>�w
�TZ�dќ��v�G�<mr�N����klv=x~��^��Ͷ����O2}$F$C������#�A�XlxVHYEB    2a14     b00�dQ�����,�Z��`9<�Ē���u��Jò��Sn��Yc�ɼ�����\غ�0�O���R�rp�y���L�YH��V�r���sv>�a�;�(mQ�pNn����z-Ȃ���H[߇�+GUO{ǋ�?,�T�(Ud}5^#C����og_$$�����JK�����;_L#ha3�:��Kp��Lm�KÎ�0���eZ(P����ʶbL��l�N���Y���|��Kq��a�<�
X�6*��8�
�-�j(���+t�y`���ok���rp�w�Ѣ��W�e��O���^]0�6���VG��s�i����7oBts��������:��!d��1����6�?�����m?����2M�<hC~�������Ve"E���2�d3U�i�K��b"@��{��=�,ڰb���eͲ�0��I�#�+�Z?��.R����@KE)h+�y�U��m�h��q1(�N:��{ӡ?Kۀ�PM�n���+�P�6�=;��K5��I�[�W�]�"}&��\���+g��Ⱥ���Ja>���%Py+������䩑��\X��3�i��0_��av����,�x���$���OR=�XE)���ՙ�9�]�Yb4>@�5�X�6��`-T8
�e@��=33�,����-�B��-�y�+e�%K���n�ݶ1aK��$2�^<��t����NuT��ڣ�Y�����@c�_
"���ڝ%v��T�� �1G�<*sD�j�┑҃�x
�lu"˜UhjV���Ҧ����ӑ�P��ؽoB�?23P�Gn���R_�U��-�rg��T8)�ρz�R�ѥN�������V:P��6\��A ���޵)0��2+X����JjIe�6K���R�&�)�M�����.g#�����&y>�`·��E�8�/^Wܿj���_@3� EH!�f,�b���L�x�s���,����;����t�p��s����[�3�Jq����H=+������F�=��M��]W*MT�ir���\=
ٝ$_Gw �T�L���}"eMY�2�tR����5i����h������S��Y-@3�A�V��D4�88��L��c��C^�R�&��"D;���SS�FYq�67$.��%�✛S���#d�� B���cF��(ǐ�s�y��!�S��4�z�\~L��,jH��*^�� o��xv�/���lO�	@t���/������$I}�A{��<��Ms��O�5�y#��G�gr�61)����;X��͏HB'�TQrӇ+2ڢ:�Xn�n�,���D��Lar�n�͢�������5���y�z����0����߉칾���[~�4�X`^��}�W�N��Y�@󓫷i'������F�<�_�P�
�������%���)�ot�A{���Y�j4��&㌟V�mu�PRTp�zx�e
�����{�-Y��˗�H�q�P��<r��f�l|��sSZ�:0�2TaO��U�C0�F�|�RWk$y:����.v?�,d����q���$�"y��h;X��l���m�·)����_Kn�2�$-.�"��?g�Qm�73����2IZ�5#(�KP	���q%C!Q�<R���q*�V�����,���06��U�J��H�!�-��=�� ԓ��v����y�a~��m�q3xl���A`��r�%��'}�A�\�6�)�ta�s�&�f�����$6G[��H�es��O`/j��TY Sb�V:䩽�_���ܷ��i#��i#¯7���4�����<�}Uܗ8�0)h�o��a&�ev�~��'�.h.��n�O㟨�@��[���%C�^-�y8Aq�$]&aR�b�w��[;��F>@��RR�`�����E8��V����=������d���O����<���=��	�Ͳ��օD��������6���ާ���9_�2FWڭ����𹂏��u<�*{�]�N���y��R�^�v135t�9(�/�ۙސ&���&7!�K@~�<<��.������74u�D���sd6��a���`j�[�/5���	�(J|�"�}%��h�h1$9-��c~YuC��:F2�_����pC}��1�"��R_n�>*&(@)q�� :GOy�9<�q���S�ǘaH>\��o�?�r��܆��Avom>�i`N�J�$hj�)���!��n�t�H����O�~��-�����@9K�V����{咵Z���ȓ�,�t�����3�$�-��d�/��6�#�ee"'r���]Ҷ�Oߏ��M�F�^��Ar�Aҗf�9���� ^���7�B.,kw$dg{2�>��M�v��XyѸ��rڔoD�|sRX�_�|u�xJY:�
�����.PeDc����X�9��x1(��>�V%����ͦ�^h���+h�z�<pj�x� �a?�:� �3-	h�]EB����e�~�<Ō�׶����l:��l\gU������5{�k�b(U��_3-e3Qb���'w��'���J�7����_�bnȢ"��	99� ��y���2;�J�o�4�3!��V<J����мF7$B}=#%|�=3'�I�}�M�Jҟ&��s�,�4+�����Y��vd@�J9���+�7o����k��J[�>ƴG�-�V�^�X���V�s�&��������.�M�ح���f��k�̦p�*ߙ�FM���������Y(�}�����O��7�E��-}�2y �� ^�7�~6��f�YǕ��2b2�H�#��X��6�b�ւ�8�A�t�Ena�C��