XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:���|�����{�C�L^D�6B�C�
=c���\6+���Ui召+3DI��~��΢�0hk�ޮk�E�����ni��[��B�ĶD�=�hQ�����-��>��P:m1uv�f�O֢r��I���%�v���|�ǊR�K˧��?�Rǎ�a��o,/�W���8�n%���^��&MW<�y�]�W�v;��C�%Cy�mD���J-M\�\��a��nd��K6�p��h+l���I8���(�4�1�2t�%C��De�aH���-@Z*�7�C��l�r�Ŕ±@���K�X�.ӑ @g?G��C�g@��ṁtʎ4�~2���5�д=9��]�U�o忡���+��.T�\���\�\d.o1�]�k����本������;��#���<>&;`͇�?�c��g{� ڞ����t� b�Cw5,pF�go���Y����-b8:HҖ�C�W���Q 	�;�H=0\��A_�q
*��R�}��X[zpK�|,}���g��Y�� ��0��5\�7N a�C������l�������/�߹�����X_���(�c�TM����Bn��g����𨍷�zX�c�ij���)@;�
����?�Lk��)�����/��.�orD����V:��B�jc�Hib�w�
hʦ	��]�\}�ݿ +��,
O����jW� /Y0�B,���'�Q��}��`��	� �ּ�H�5�1��
���c\9rz�n�*XlxVHYEB    1f41     990"�� �~�O����</�
�s��<�S�A�lpܢ2�]*I����g��3�J}r���m;�^y��	��d\�c��f/Ӗ{���~=�{��%O�:X"���֧)�jʾ�i�9�9����&#�o�gF�^A/����C��:��s=������P�P��}�ҘyH�3KK�
�6N�0Ý� R�4{OJ�Ne��e׳���9F�T����$��Y�C�9W]�[��TxӺ乿Z�>=l���c��Ï1������I�ʯ����7&}��`���t�|���;;�Q�fv�+����;f���Y��{^�'o�O�����&)��m��V6I�l?Ժ���zj������|�P-�}Rq�SW��_@���&Iնٲ�+�hXb��˿�[�H�:$�\�vqWK��"���1�J�@r9$Д"����|;ix+��[�N�Wy��+�@1��|�Y���SX�$.�S'q��0��Q��v��Y�pXRT��D�q����eb�A6��J�បxau��
2�=��zX�j����n��T�X������*N��%�9F����t0W���T�߫m��E�zv�y=�O�L�����H�.ۇQ��w1��bU1	�\��<G�P�qEG&	��)�P]&r������>��b�����W�v��N���y��X��҃#"��rQYN�?C��������ξ-�G���0�>�(��߬S^b;+R�/�)R�4�@�dõ��`�5��j�*7\-٣�Ю
ȿ(�_���^^)���km�w!�΋���?_s����)~Ӻ�;��u���C$��l�� �~�w�JE�#\�� ���!x�6k��~!�)^��6��i��U����hhlV��_�I=�WJA���+X������$d�ļh�H�˺����nf��=�l�Ŷ���6���� [��\d�c�� 	Gh�ɹ�3�����aQ��}RW�Z��C�YE�4	޵��QU���"m��xT�{<��w'�U�c���D�g�A�
�i�$���"�8���O�Am�E�a���/B"���`����kd~�u6U��_N���a3��W1��)7V�x��M����^���t
��Ԑf��¸=����E��*e|E��%�޶A'w9q�@@D��_���W���B�͆�Z��>�tT�ł��9�V髂��7h?yM�]F�бM���U���L��2ĸ��Z��{u@R&����T `?[�Ч]��
�4�O��<&��$-;o��\ߧɒt������d����^�nQ��~��p�!8�h��s��fu��G��"`D���{�,�
��� �sv�Gq��*QӈV�"v��?����J���h��<}��`�4g2.[gb��=0?w�\�|�x�ī��͍���9!��u`m�����z-��+�>��gBQ���� ��(�)��**���`S{�SW���۷�����U���#�OJ���O����zV��Q	5����\Ԟ��R��W�gN����T�I@R�$Gݽ� 5�9��l��dw��Œש����Aoh��_���&r`A$C���<�b�)<>�_m�V��k����-ĩ'�L��9�Y5"ñ-�҆W��������U�"�J���4�k�ǡv��W4���(> �"?��~�.�7�Lu�^@)�����xhZW�dʹo+&����l�"��k*���g)����j���;V�5��7X��|6!�1Cv��,G�O�g��w�)ʫs��P��69 �dQ���2�`i��y^��`ug���|j�u��Qsi�69�?�ɻ�F�E��ȏf/�֫kwױ�J7fe=�{������C���ip���^���	���5{LKl�O��f�^ZwC0O�S�R�C����Ҟ��y^��4X�M�p��3�j�r�"a;�v>K�h��ɓ�����vY���f�3
D�уh(9k�nr�%@W�Oz���J�>�/BN����~:��������S�pS�C�ԫx�L]Ď����ߪj~?&ʶ�g��sieٳ̓�@���:n���K����^�C�뿌����{��2��b�@�i�0c�1��M���J�P��L1*����c���"��*� GL0��-������oXlℨ��nx�����djϬÊ&~����ڥNV�0��/!t�D ��n��v�~1Z�	� �W�Y��P�gj�m���3B�q���9���;k�IJ=o��R��n��4dT�:`]b�M�a���oD������
���ӿ�V�񱙵���\�׏�ɦ��g��lu*��%�s��D��eՊ�s䁩ó���2;"A��!���a�vC���j�XG3c�� ����Փ\��m5/+!�M�ϣx
[|<���?�Dhg���wg�Ci ��DV���
���0�>n%