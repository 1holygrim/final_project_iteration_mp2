XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J�\G����7�D��.a`��j7z� �.�Aq��P-���5���S��k�W5��L���Z;�]��[�X�B�^"�Gy0d���V~uF����S�Q�ʭ^ aU��k����{TS2�q�߷�1&�8�T�������!bhCb�P�O�~Ef��@^�]i2ÒJu���e9;\O.�z��W��s$Y]M�[�+kWP1Q̍�����W]S|=�^�?&/qjg�YN|�Lϔ����tL�	��lmaRnh��]UW8ˁ�Wyd�p�Ği�8>�h��L�T�.چI�/8��Q�3{�M�%`F�������vrIp1�U�dB,fc�J��%���Pd%Z��65v�knZ�H�2��:�hK+�
N�Y�)�EFB��`���!�����V�2I�t����P_��0{�R~�LU��M�M	�S
R�]�m���-)��Ʈ�9�F$�iB[0�ҝ7)��Ԛ�T~3O&�v�`���1ly�
�-.(�m��_z��K���(����bWtF�K˵�7��:�Cۻ$q����N����*��:6~>�mL���jM�����θ�M�{	B��5:��ڱ��6~h/�Ԋ�z����;%�xǾ�jx�X8ÛH��%'9����xe�U]P��}s 鮈y3�Gwӎ���_����I��!+K0�G赺3�i5�[����Uo,��x�Ȅ����=�Ryo���iF��1���g��%ۮG�����XB��a���!��1J�C���XlxVHYEB    b087    2540&�OE}��ϯ��Cޞ���N���n�g��i%V�/�K�m��*ԯuL܄��	�9�B�j��+TMoyח�	w��n�M+���I��!Vϕ�=ݖ��U������-�WQ"oI��i�M@+�ӗ��2�@2l�V�/��I$Ӕ�5>��u\ylG)Q��}��K�=�A$��@nsQh�3���
�ܝqg�i�T�C�_������_<]?vH�WK2��.C0�̈́ՈSGg�ڌůb�v������`Y�R�f�Ď��`to��#o��W��
T(]ޜ|D��Ƕk�a/�є�4�C� ��>��l�՚,_>V�{1H�<�$�W���(db�x���˰?�����E_�l�`BLNϊ��0�\�} z;w�O}p����L_�xٔ����S���=*�����#�M�rG��$LY��N��y�'f��ݒ��_�c0wW��=���8=u�]�T�����dp�S'�~��$�@kn,pQ��ÍAS)�8��x�	�j]�Z��PK&�t��&�\�}�h�ӷ�5<WG��bl�L�v-�5m��Sq��S�	ّ�U�5a �Ƣ���KS~g�h��;x����� �vW�ٌ��,�s�tz��h�� nH�7m��CX���czVT XN�ؠ��΂���V��S��ho~���H�$a <�8}�8F��ƿd�~.	���hsY;<ss�H*�|�Apw���r���"����?.=��ѥ����hIn֭� �H���7���j�#�sސ�����^=����;��T��/�l}����	jGt���<����W���!�j���b��Uz���$�2Rϫ�V�4󆽴�v��'��=�i�*)̽Y^І���yA���@�L��*�]��)��y�d��#�'{�4�C-\ޚ���f�ߖ5�?�ܞ`������f����Oc�T]2୳<�cu�pk�ix؁�lN��\�jr �>6,�:ad�e|���n�&��O �C��6�a#X�!�:���^���x�U��@0�r�]7�Z����^�v�nF������fL�R�"b�h��q�C��N�_�?FP<Jՠ�@ΰB�u�ݬ��z�8/�=��u }ӷg���l�v��^��ID�-_�ǡ���F� 6�8=�k��JJϙt��=�88�����Yϋ��^�m�54�7�u��w�L�Q	�������,c��5���3f%�q�(�M��0��:e����(x�V�H���!�]�H՘ސ��6��Ŗ���k��_��&���pgĜ���y`f��xw�s�:�4RM|$H�uM]�Bx��P�8����4�1��o����!TP�t�=0DsB��6j��+N�k?w�
'%�u�h`&�2���65�WG�5@������-�g�5/\;`�l�j��Չ��o*��E-_�<y1�V�w�dn�GeH{4; �nρ�'��.���6�-Iz{Pk�����.�H�5���.�N;��K��<H}8y����k�e,����tϓ`6O�	]�¨Jf �6��Y��B�wR�'��ɧ^\� Q�G��ۛ��V�*�j.�GPo�*V����3��S�L �>!��>J�^+��1{%� �qW�=�(m���Z�������]���Jh&��픘���e��M�R�B��{��~sTtŝA��>�y�S��mW��'����	b��LICw@HRA%�q� �����D�
��Kʿ������M�'�|k�B��ʿYcL��(�/XX��l���۽�)znp����E=�Z���f´��qQ%v��?o��k�x*��O��r����������u*抓�ɗp��bи`�姓o1�11��>���(sԂ�dkayc#�H�6��M������M�c4�cṮ��͆���>Hx�Ñte�jGn��M/+#7Bd��@�r�L���[��9T���ky-��(u����>�=E˲&	y�$�"/58���!TQ��<񛿹���� /M�Mt5;����U��b90�N,�G҅?}j�є���bG�мopȳ�%������c��c���Յ��7��sQ�0�|��e�Q���M80HƟ��ɠ�ܿ��nU���*���y5愅�������xd��V�3���l���1aW����o=װO�2y[�Xpɹ�;xӦ�������|Yc����C�Y���;�+LȦ�4(s0Ά���E�J����k�6�i�ȷY�7���9�.�D�\Ř�������}h��8�[�k��E��!�?�}���
ٺ�c����a9�#�a��d�CW2�Μ�r1�ڰ`��.R��S3���׶�������p��!��[�~{�5կF��"KI�`Э�PY�m�k>2?a6G(_�W��W���e{b�}kCh�7(�%K.[�ԓ�B���iӜǩ�I`�zC�����%�9��s&�
����]���8�y���tTѬ/yO���̌����&H�gB�d��f)�Gͻ�ݦg҂�?q���>FpG��]��Mx�� �$�T��z/��jQk��)�ݝ����|���T�'�.N�i�_QǷ�x��.|�C���"V���u�s�)��PJ���2�� (Gw�>w�}��@]��A�U/H�jڀ.��"����k�M/T��ܸ�R��� 	.�7ɞ��u�M���/l1��$�"V��	��[8�&(g�)ǽ	��������&~]�i3��ʒ��� ��[��YN�V���>�
C�Q��i�*��M���!0x�ux���_Z�'t�@�d>�LS@�-V�irAe�y9�Ta��oM�M_�5����7�W,;�Z��tPy%��c�����B�m�w;^l�p����[S�m���D�4�(?��+�9��2��"��.��
�Ϟj���,i���@u��?���L�V/^҉T�JF����C����ګ���c�G���Ĥ�{��=�2Ju��`j:�OR;W�uG�ȟ�Q1LY�M�^4���N75ڊ�ѡzf�"/��Ъ�QR#�I窱�I�b2�yC#.��� B3,����A��ڬǄz�_K���^+T�����Ǘ���ԯ3"�>Ǽ�XFˢ���)���8�K���NkCt~C{Jie����>�K�D<��L2$(�'	�_��gܵL�<K�,`��c���H�$�}S|�˔ݹ�6����Њ$៺� /��wZПݚkX^���h���2LµP����Ӌk��a�K�|b�w��3(������Ub�2��	�����o��@��Hs�)X�5�$�L�^}���Q"}kJ�}T�@r��S<�R.Y�'B��G��?� �pww"���y>��?X8H�lQM�+�p^���~�F>
ia��=�Q��7�"�P��/
���o�y�#�,����[l�h�I��#�8�oA8���M_��9�9Ȱ�)����.sZ����%���Y�	��AX�A�Ո���l��"ALRP�.ʁ�G�f�ч�Z����f$��6��F��F��֘���ɏ���w"������*��4 U�sl�k�ⴊ��k_��HrϾ��&�e�3�yZ[T��Ĝi�5v�k��}�����c<����eʎP{V����O�E�l�n���e��P��-��Ǎ	�s��V�y�B�c��P�Sxx�����(>�,%G#��?b�ÓOu�{����R�E�"T�u�
&�\��'��-ސw&4�X���v�Wʽg����$R����;�g]��C�ܙ�8.�v8��M������ĉsC�pk�*ĺz���G��vt��]�# �b��d��~'q{d9��v�*�<�g�OL�"�!��99��p�r��1s5�d�M6&�W��@c������<] �ژ�\��w��N�ΰ��)��_>�/M�
����2���:#�į6,P�غ׈��7�4�_��S��ʪ���z�p�C� ��:U�d��z���;:��7�ݏ�I@��ec�6���W��6E��ۮ��\�����E�:h�袡^�T�\�}w^��0�G;,b�f�5z���%�]`���1�I8�]�±P�y3�'E�� �g'�#I�u������`��.X��ȷMU�|G��[���<�v8�~�����E˘��3�Bg:H��L�����ҢF 	m^�����2k�yo�=�H�>����m���S�9�2��"M�C(�c>iDF*�`զJLcC����|gp"��o�xK9X�Z�q�q~O
Ж�U%��4NO����w����{<�1��$qY�^��3{h��f�rI�Ȟ!���kpn����s=���9<�b�g�pb}�H��]^�ᐃ݈���rf��0�$Gٜ�<� }�&WӠ�W�z�&���rgt�^��Ӟ�y@-���)��\�N�ޡ�L !-d��ր��a��_���T�hT�R���Z�unf��AνXvˣ���d	���iGwVO֊~!�^h���[�k%�uK�~�<��ĭ
���c)u��j;A��:U`��[ܲ�;�[#yI&���F'���И6�-)"�S� r����B��k��M�ǩ�����P��!P�#��_�!\������"tB\�(s�MhuӞ�y+���
B�=0�A�/F3���ʤ^k�k:J����������^���bt���@��4Zr=U�,q��yܑ�K~h��E쨆���q�4A����U���%]U�WpZk�M[~�����6f�=y��5�E���}�u��J�.If�Ҹ�A�	U{��hE�]��e��PzP�h[l���9��'���\e��S�����57�{�M����g�* ^0�Ό����^ú^����K��yQm�m�)g�a������zQ�3�a�vM
���a�R Y墾2������\��ȅ?�$v�{v����o��+������B'G]�H�Ԑ'�����_�LuQY�F21��q�^�	`N� LD�n�4p�O��)')�x����K�Q���^���������v޹����6x�t��D~9%��~��a�n��!t�Q����H=B���B�v�mVI;Z�u�2s��ay|]�F��lc��5�bp��O��q��!Ն���S�,fy���AG��ko%���ʓ�YZ���S�K� CR�^�������+ �@{Zy�¼s8�^��vh�K|�р��a����<��txlư"�DЫ�g~��t����暹�BE��"t��Ɗ�k �\�
2��C!�/�����b5�V �M�#����8�=�.���  /�� A��=���/���G;�{�0]�'`��>�������#N'��t4���s�{�Z��;��n�>�j1]�ɔ��!�
��j��&u��q�|� 	A�&���7K��dv�Ij��B����bԁ��x0� ?��x�\j�����Y� ���޼��X\�T!6+�\@��"�<���rH�$5���������� �	-������o�rz��4x�X��hfE��M #~�pEv�򁱇M�`� �h��}�� LずӶH3�a]-�D@�B��5�I`[W�#Gd����x�5}�\"|7w���i��xc�/6�Ŵ`�W��0�E��k�/H*��cU�Wk!wI�k�����υ)X1�{?^$�/@XZ�u�ή2C���nD?�����������N[dy�Վ\|�-��_��zy��;63���ڨ�?�\����UJ��WY�^\#�$�\���i~����9װ*�0>M�r)�#d���8�1kIR͸��������2i�W8f�`Ȟn㺝�!A��e�0"�4�n)���O�9rT|��z�������.�&9Z���u��{{�e3j@��`̟Z�0�"�u����x��g2 �C�D�����gC��	)��!P���»����a�EF���_�;�+��)P�m\b��Tٺ]G���6})X��j�����nn�M?�k���j��"o	�����ۈ�H���	Һ�7QC�ަ��{S��*{y�꒝<�K�ǜIOO�=�r$vsf���
�1}�z/�?y�G�C�G��ܰ(��v<-X[?y��?��Ƃ�ZjO�8����6��>�g����r��l*!pd#��%|�ߨ����*9K�����S��#"�!kO����l���, *٥�&/Ү"/@ �r9�M;A�cr���@�כ�с~H�0S�(?J�'���[�L���o�P�����@�1G|C@<��h��UJ�|�x��%l�RǝA���z�wodW��7J_BT���!	�����6h��a�l�� <�o��N+���p��V4����*v���P�f��.h��ZGMC��(4h߹EoG�p]��ú�5G�~t੥��z,OK7�ZT�l���e�+����( z��m��0-Y�=&��bt��Z�}�G�bAZʅ�oP+[�������d"w�p}Ro��ٖ~��rAOc��1U6fm��>�t��U�"x�z�AS~s������Z>�깫�T�cD�#YB���.�;��rxE4�YOV���g�A��#r��ƪm�~�/a;�����n�Û�M�t_�Z��AI���cR{\K�F�&p��o�dR'7�)㑎&IzN���N�`K���1^f�A�o������/6[<	��{���ǅ��|Y"˷v 
5�V)	7�o��7&q�!���9���2L(�����8��lhn{>@���e��3�jg{,���x��-������� �����9\g���l��j+��U(�b悖e�^���o������;��r�/L�@�85��L�};%7��Vsrc���U�&��yd�}��UE~��W���7���
JXk�Ź����j#�:�S���v�몟�6����nc���1�cU*��%����u���m�;��<�w��8%ć�	Ԛ�8J��\8o�L�f�7&ƾ������.�Ʒߌ����_8�OH���ƍ�br��L�󧉄�T:'ş���|��5e>��W�eu�F�"=�y���g�˷㠗6��>@�U���>���l�Th�[�fQGy<꒥�P�Q�����4��b�*��BA��~�D�g)�G���UN����o=�������gZ�=S^x����jc���Dmc����7�%���r�G&f�(���F�h��V�ӹ��b�0� ��sr0rZ�������Gk��RLg	��7p�0� [���t823�}/Q��L�q����r�lWhہ��H9|�Q�Ⴁi=7%�}&-�("�X�g0n�������펒#^
%+�q��J�Z��̑
�i�d�:�\K�5)H�r�LЩ��2y���庐 Y�g�^�q�����TH��$<��]�5���� �8'����Lj)�cuz�v��� �G�����e>�O�c���ɺm[�J%x���/4���0ŷռ�/��O]xI3�҈FV�ɻ���\��;H ��O�U
Ş��0��d?�H���i�	�0�$�<�%�b�g�TS4��qД�G���b#�)�dN��gcd��2��d)폤Ҋ�R�%�e29 �B�!����X/b_GB���M)ԏx�5ir�ĩ�5%�v���]� 0����Ju"s��^��L���ݴm�@��7����@�ql��t'���
;�<���c!��w(T�,i��ā���c�lY�Ȼ�V(T7R��"Q��.X}�}�5��?)��f�J3����@٢!��Z	��t�r �a2�Q��j�3y����O����Iy5�s9�g��P�~�Ss��HS�;�}���p��ú@$?��@.�A�C����.��ZQ&R�6$�@��"�����A~�cڌ�8�����W:�Z�3Q솀����
}���j����Ub�PÅA�Հ��5�G�%��#?�3��~��U��t蘥}���XD�T�y�ʗ쬷�ڕ��N]G�͓�s�	�i5�HZi=\�+Q�Dy�B�-�:�=<l��j����p�U�L�Dg�ݟ���|m��p?(=[��*D�sg@�C���.��y_�g��
5��A�Ȓ��Pw����uB��3��7�kJ�J�z��5K����L�Gɷ@@h�"�*���L��3�_��v�E�#�k-��V	�@����%�Egw6�f�*!�oHy�TƊ��η
0��>�v7�/�~8z����]Z�y���yF�8K�h�Z6=�(G= �S��2�l
�5��)��	ȸe��k�H�����Ԋ��XO��τ6)F�������LVZƢRYsԴ�Jv�S(6_�B�G�W�k;(�Y�^{���F R��A�B��Mε�.
Я���P�>`��Z�9����]��2�9�s��d��n���.� `c�%�E(In�&=�)��3b���:�����@n�s�(	s�3L�k�k��&7��cq�	���an��B|n��8�kz�i���f�.v���#]�N�;��ǎ������-7�{�DmcO�
�s4��L�#"�)��Ik�h���{�V`�R���B�0`Kzȷ|՞�hs2C���AP�bOޛ���`����}�~� �4ˇ��MT��r�c��˦L��R�hN〘�PŮ~�3��!��z9� � ��,z�@��D4��V���c�w�(Zh�q�F^�g��RB��+d3>�|�U����D;���;Є�b�����I��2ֳ׆I��C�K�%���\���W�"�>��Z�,�L���3�;賞�
{N�vf؂h�Tb����E��jV���jn���P�t#��C�� =y�@��o��w�0�<�z�/vjW���'���#�3�Ά(f�Nj��A3��"�+ë��R�Y��|��"M�"=L7@��n�	+$�|��WX!F�0��ＰK=۟�����kta˂�3�@8�Hͧca���N���1.ґ�s4JJi�����յ<bӰh|�Y������Jӑ��3-vRJ����1�0Q�n��o�ʢt� /�v����t�ɷ��
�-i0K�0De~��|�az34 �I(�_z8a��a�n5�Y�h@��C�%z	h�� �Ϳ2����L�+���M�3LG�p;o�P���}�8 eX����bc�`U|����09S���)�J�*Z�H<���'�lV_I�5A���������W1}$���/�Q���)Yy���s�K�l��`"��@gB�|ֳ� ��@M<0�ma��z�g��#���8R!�ɠJ�����.h*y����~,ې��o�M��w��Rd�.�����/3MN��"3Y�XMqNޞb'�tn����<�1W(}�6I��f�P_mR��+���D��G��ԚM]��O�@|�a�	(�w�C6Cߣm��s}���=��\��^ʜ�"{�'�`��cؗM~�����oi� ��� F��N���P ����}|�P��H���