XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&������>�'w���7�ۼ�0v��.�sӹ�5�X���#�)a���\E֏����L��W= ��O=��|>��(*#aǼl���]rk�`�z�K��������E�!�S��F�O�9�8U�y����⽱�<$�U�
�5��v��Vĕ�Vy'=~Ea5���l��Ox��>cH��ֱk��2�[��Jx�g �K/ �6�ۑ5�䀀�waM�_��������+�	�kJ�~�c�#�i���{���^V�4$�m�36^S_(0�Ma�ɀ���0����2)�o>
n��U��
f���I��c=�c��v����5������ xf.������f�Տƀ[7b=����@�P,{�S�ڃ.�AX�1ʰU�P���������V�Y��؞^y;k3F2m�H�oW�E[b��km%L�yx3���p���~/[���2a��T�aq0ǺZ���@��Q3�;SN_x�l+{��.ѕ6O`D`�n��"��Z\�`����!�u��*�	12�袅�&	�����-�����D܌ɠ�*�I ����%�a0)o�nC%��%[����$��n�f��g�7~ɼ�[�J<����d�n�k��J{���O;$
o�\N3��Ƭ�Wɪ��G_Exx�}[�͋�T�h{ �]ZtT����F"tC�۝!T�2p	�͟r<�]&��R�����眀o�%X��z�3�(�'A��\ņ;UC^��a9���Ƭ�����o�R��5XlxVHYEB    30cb     bc0�������| b��3?�����mqh�K6�[���s,���5��J��,-�G��P�ѽC�D��y����Uh�Q�����ɴ�c�w�XI.�(޴��yëN{�-�T{�Xϳ��y��㐆6Ee��k�M>��}K;�&q���|YO��f1�:��QΫ���Ȩ�^�;rhT��&϶��Y�å���6t�s�� ��f^���rV-1��,)gԏJ3/��"�6��69���}�L����9zb��j5c,9
؉�˺��u���V�O!������d�.���\�ӀJ��J�ۦ��@:�eVzZi:SN W~�PLb����v�<bv>��|u�\Kt����=�J2KRl./��^��P�/�c��@5md���YX���1�;���/�(4�\߷Yb�'���X1�@\4���F������ؿt�\݊`���aM��F�ؒ ߞs��ֲ�:^$��&r1�-��1i�Op��C��d�e�4��̤ �I~�@�O���	��Pޞ�ԋ�Lq���dr�[��]{IZ�V�^��Y)���Y_��5������)v��u�.A���-�(o�pz��v��v�����7 �i �!;q���#�2�kR#��&�8����T<k�ɥl"8��O�~]N�q�)�P�ss�I+�Z�$/�aƗ�����42e�ٖ����(BLU�e](p��=i).~~��Ns���6R
ZR�3�+w��.����M³�[U����`%
w���	C��<˂�>���&�A"\ф��~�睋�9�y6��19 x��D�e����U���QA��	^�_�s#}�	k�Tqk�5$�k�Zo$Y
�=1�T�ʤɡ��C�A�s"�������y˱����Fo�����4۬z���8�͜�A��� ��9�/��P�:��P���S�A��TV(+_��ᎌPÿ"t �7Y����Ϙ���yxR���H���h�[������)���Dʜ���S]Ҍ<̅Y)��Y���{�M҈2YgSXL_����$W8\�̅UXZ�`�h��,��Y9����,���rx�X�s�9%�t7�o'�|�,������vOQs�'��kh��6�;��
���r�V�^���.�����Ļ��jձ[�i��V��]�9���^����h��O��I>)F.\?²r�v["�8�>{G]���g���d���4u�������GmE)E�qe�R�I�_��gN���;�.9�!���:�G�ݿI��	�K�<�,�Xf�p0��1���.��b��j���D<��p|�@�C�f9�t2����}�w��ʩ�_�e�J�Lݳ�)�����%A1�����"�wqR�`S��L m!�Bl�*?�+��ދ��R�%�4�U����
�h�$5p=d;��FK%1���3���/i�I������];���!�E/� t��ė�C+�qZ�#w���hЁ~�)7�G�@7g��
�_f���հ1��h�y�%u7��&�b���>���G��h3w,���7�b�I^�ǟ^�aCE�@�a�u��~��eF����D�h���4 _��o��u��5(�b�w����|�1��aj�)'pƠ�A����U�9Q�$T�����M��YR#�(~ 驯Yr��þ���ժ�q�Ku)�
���)=M/ Z��μ�R����Z����>q�*Dgnr~N�BwG�d��`	5�5�X�تg����c�A.F�'���9=P��j�Q������W���,
��k���HSa)��d��� ;����j#�;o�p��xNX�N}5�m��JY�_���m��g{^J��I��yҦ�Xp>0ML��i*�yq_>N �<��N��5L:�Gê?=9��E��3���t؊�bI��U�n�����`1h5�I�:�fI�����'*1΢�E��%�M���k��OtR�7����}��[�>>�;m��g�����	c�h��(Οn�/��:Nj�u9K*@W
���S	��A�<,�"eZ�*g�*���#W�������z�Oh�۽���?���*��h5���`4Ec��螠��D����k�0��i��3�YKc�E�|u�ӌc��#�2b�h(�(_l8���w[��G��%aahG�OsOF(�������"��3aȬ���e�5�fx�,Ğ/���k����g�	̰�wSH`�\��E��5F���X�xJ��(�U�9n�׻x�
���-�_����F��;�����Bg
6�5+����e��x�̱|���c����/�J�Ç~E9JO'�M6v��4Lf��u��܃�z6r�V2ah)r�IB�Y�%Qٚ� 9�gW�8�H�rJ���E�ϗ�hBg�-b�����YM�d������oR����V�O��n�Iy���_�%L�R�;����=�.]	s�d]B`N��z�k��s�< O�'�F��d>�+O4Rjd{�gT�����՗`H
��כ��C�5�0n�Y[��s%eKu鷠J�Cld�T�/���q�M�A�1I���?l�t��R������a(rk�z�qe�K?C��)R�VJM�n^�8���� �� �O���ߘ�9B��v��"zV����t��{�Oe �Ba�MF��X��pHh�����z]J/L�[�#G�Zy>����Ta�S�{�7�!k-.�1��>�u��Z��p*�I&i�+������nŚ�ٮY��ll��J��M���g�%�YC�S�k��A�׋w<q��<�;�>�)Hp�> ���|c�Ε��,���"�Ć3�@�wa���Cb�H'G-us)	Wb�@�y��+C�8��J©U���Ь�P�c���v�տ�h���uEH:d�a/JtƍG���|��d-
_��
����(؝K~��s|�gM_�0�2�]Ou���X���� ��{&���	�<�0z{���:hG