XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���,U��VÃD�y�V�i��'�N5�4F�:�s��Xv�)�x�n]
p����J�:�t��[%Ҫ�>W8��3gs��0^N�/E8���K�z���p�tWT�.���-�[�j��r�{BZN�|�OT%1���Ŏp�jl�X"_��v{U΁F<��������X0����{F^�]�z��C��]i=���Г$�_w��Vr���, ���(hd�Ӗ��1�C�?N�D�f��9O"�6YI��[GE_i�O�{��{)�Q/�����.z�̒M����-�b&���X}�y�ڴf���~�℆5\��*����S�S���"�l�I��q���@5i����'8�1D�#Q��P���f��S}�Sc�к���wր��Ff��υ��r�񱬻:]��2��r����*0(������I�͈�"������A�TH2E=��̩��H�k���.�UaWY=��<��KCT91�&L��
�؆ev��ץ���qԨBg�ս��t�
�"����h��uuǂ���Sd����8�R4t΁G.��G��V�Io�/����_�N����xtv"ֹ�ν�m�2�������1�`��R3��Օ`�P'��B��t1΂�x��x���}�>�`�T>���~���l�x5W��]:%9}��f9Og��x��R�20�1��.EVć�^�|G�šģю�-}fO�r9S�{�R^�SݷLZ�ǀgr)�x�i��("ߒ>Ǟ���"��N��	eU1�XlxVHYEB    1a0f     9a0}�N޺T�U��W+�&�.����=V�����"?�
�����f����_������u9�#���s/��uo��}���GIm=|<<��-GU��IֻX7�ߣ✪_xSk'��`�!Dj5��||^�b5���̡�֒׸�Pi��������g�?M�*|ӥ�Ņ%z�h��R�k��q��ֿo���g_ADa�^��
t� ��]�3��S����r�̓s�j��
G�r�1�.��y�⛗W9D��L4e�C����۲՞z���gc�Y��w��_����=��h4��w���k��zr�xj-1�m)��H��>v���
�X!L:��b/�����`ܙ�Wx���Q&��մ��a3��+�-8��f"�N���J3wy�!s��.�͡��A?�Xv�1��TN��B4.�^�2dq�U�:�l�B�	e�p��Xg���Y�7��FzT�y\��NE�Pi�G4:2J���U�Xb��V�J�e�C%�v8iՆ�G0�Ә�1@�X�-#�T$:u6�b۵�3�T�<y/�0tI�1�WYvk�o#�[qQ�l�Kz��ds�1�]��*㸒;���|���j�*�H:v�<�}��}�0ޱ���E������Y {F�5(C�93�ea)}��ēb�J�7zs8��=�#ƄvR#t�n�PL{y�����d2�Մ�07�mR��X��&�FHp!3}��H�L=�!��V�Xs��bzH��	^�XxǺ�W��;Ʌ-�4�kp|��g��θ^�+��\��J���'7~�R����P=�i2����x�8#��*�-4�Ź��/�j�p�,�7Ȩ����(�/`��kv|����t.���`8䆐�P���Y�B���4���ۀiU�ԟ�V@�Uo���W�f4)��h��c�_����DP��Y���M#��x�u[�2�+U�N�y��Ԩ<p2����e����q�R�ebO�T���"�[��Ax>��� ��z@��&�� #����������ҧ����w��ˢ�%w�W�-��	�e�	�2�X�7x�}��
��t�4_�F�1k��sW��R��5�F�K�ا->�����jvWe^u�)q��!poc.�_�����SL�i _��Ԏ�1L�Ю��ajnf�ʹ����<|����C[}�D�b�{�~��y�tq��Sq�#� )�4�R�[�4����W�� ��/���:��$ʏ�Q��]z�м�җ`N�c�w��	PA/&BH�tǣ�d���ι-!��r�H��-�\�c����X�ڝ&�WW)�.q|�]��m��7���]-	kǒ~>f��Š��~�UZm�fKކ��ʭ�X�*�э�/�F{SL-�>�T�4Eb+�H��C�-<U�~����u�P:e*u[-��B�G@��.ãlT����@@�Y�?���Pf����RDX:�
#v�#Ƴ��	0>}�?��!�&�6WA@"p�6�$� ����"�=��E�^�gƩ���ԅc�^�^!��<>��~��V"�pݹ�=���?̶/2��RH�W=!G��ye��������5��`��������`�7|�Ц,���Y<$kB�2��7�A���f��Ky#��-N��%.�h?�@J��'�ޮW�M~�Ofƒ;��oLe^��B.��2xxr��}ޔ��]n�S-�	��͟�3��"~؂���N��P�}�u��XXj�q�n��P�;SA66r��y`���#�o������ʡ'��c};�Y��(�}\�}G�ӱ�x4M%'h��3�لC����μ�����R���!?� ���+�9�J�d�jZ������v��J��?������x�� �Z�9'��-WW]��[e��E��z<�ý��(.����C��j�/�N���F���O#*CV�T%�<3�ȗ:R�~jz9�/'"HZ��Ф���".<	̾�D�Ũ��e)=
 ��~ ���@�";8���8�Ĉ����ra��Dkh�%hG�����f�i{��&�/��^׻zB�sX��T	�6^Ð���YV$�Q<dI��
 ���V�&��DMu.;,H�G�%���	�n���>P��#��@`L�T1��>
d9D$ *[t�yK~��P_u,�n�!g��`4���c��*��J&�'�K��	Fm#I�U�����yNL�մ���tb�$�gc�vCLY���)��?2�^�f̎up��Y�v�ްJV��i���f�L��a`�X"��sT�I��"�OucUY_pI�����DH~�f`�&nք-�KC��
e��\�;@Xf��1�
�d�XG�����p��2qv�ho�ҟ��.I	�P0`5��2Ʊ���8*��?�X涵6�&f^땰c�#/9)�p5gI(��Bj_l���>I	%��:lP�a��8�N�_(_�n6�n�=Y��K