XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z?��V�bN��3�˲�c�P@�@�/�Sw��8J0��L
����|���K(ʶ_�]	Hܹ�)����`�m�\�A0�����R����N
��oj�����#����=�3���,����'��, z�X"��@Hݗ�yO��c�.�וӃ���()�9��9^+�o��Zb R|{9�G�8-O�o��q����9��m�A����*�(�X��7"�3�~XY��X��ȭ�D��ߠ�������\�vAG����e&��>��	��l��Oa1��h�֟�������RStu���� c�(��ח/��^O���7��<��h����w1�ެN�w��gc=o��h:f�*0�."�LBe��to�17��1KYWπ��ET��w�4⺞�N�����!ɘ���$�+�m��>�����j��DG+J#���:�|;�H��j&a?�N�����w�	Ka��H���ځ�|�.v�>e�7�#?(�=���GQVs�M�x���P���A6���6�d���M7����z�/�!S꒬�	y<&�����~Ȣt*c��E�^:O�`z}+b�"TpK��/��FeLk@*~Ө�O�-��HC�<�q�� Z�Uw��W�4�pʗ���9�<@B?�o %�-�%{}��2g������Y^���*$��69J���V@8�)�r|Yi����+S;ڊJkC����{������#�O�W�����G9��#ӂ�z]��ȹ���8�0��[*G�3�n��-���L��XlxVHYEB    3fdc    1160��C�/8�RV"���[����a�Z����((CE�Z/~9������W�ݷT��q����wQ��鴹-�M�qf�B*17����)#^n,����=_�� nB����l��{C�iǜ;�v2��Lzܑ)w�:��q2jM��e��E�q tB��rm+�O�,�\C�/Hq|a%����ʇ���%����/q�R�GU�X�&�'�-ab^�5�:��C.�"s���'?oj}53�D6� Efm���������'��y�`���������@o��Q��Q�<4β��!xf��3h�ρ�[�d+��$L3Y�2ŵcƊ:̄����ճ�;�����zO��m`�'OG�$Ko�A���G���`��%etm?�8�����8��=�e�G�E�b:vT�Z��U���<=����o��D{?�Y*�$�T�~�2M, V�?xjB@#�((9Kd^�,�ֱM8�;A����cС~`�(P��2I:M>�"��y�ݖ'�?+Q����C��9%{�eg�ӑ)��*nM���O9�W#~g��#��n��k���f?de�;�6�t�Bt��-��}�o�g�Y��
h�L&9\.�}V�i���*��!qçyLH�p���K���xv�&�I��.{��]����Wytd�fCu�J�
%�c���r��fJ<��C�Ệ2�mX�w '��vذ��􏆅h���%*6D�m��L+�ڌ-�	�n�7����Kj]������ ��L�|��]������Zi"��Tg���I���
�o1}�ӣ�۳O��~��#���W�����;N��5�P�=��O�A�����������NA벪S�Y�t*�wr/q5�e��iv1K��G�`o��ȷV�ſ��_��W7QE�:6V_��%P�n��������!=0�5�f���Je�u�yo7�7�Z�!�M��N��$��zpZ�e�}���(h�ʨ�s|��'(� ��غ�Zb�@�"A��W�������O��(����&]B%��� �,4`�Q��U;�s��h�L�%����UN!�Ol��7g���F���8vP��ln;��b�c�Zu8��
���W�g�e��♗�,l�~[v؍�r��,L���B��KO�k)�R�_M�}Q�kň��f��G�J�m+.�E�d)�X��"k}�h�!��Nv�<�(���!�?� �*M�0��[u�6�Ox���M�X��T� }��.����|��Ek��^��rJK��0��
S_�G��Nid��f�?��gi�����`VPF��NI)���y<����|[�j svጆF}�@p���K	Δ������AO�52T���(.`	���R>��ш��m��c�m����Ʃ���\�~��94NAZ�qe�؍YV�#1��H��ZØxE��z����@�IW1<�
q�L�iTq���jRS�`�������*�2�-���_�¤v��!��'�v�H�o�!/u��r�K�1¶5�\h
��u����Qj.��������ُ9�d��Mb�X�_��19�3C�c��?4�a���xa
����w��8ǣ������ �D�k��_:�r�(�٪P��̭�GG�WH��>+�0D<�A��i+��X��uP�ѩ:6��!ߤD]T[�Q��ЙU�Һ�6��G���S��q�^�`Q	�N��e������C;��ndr��� ,�:I� ��C]Jݔ�[�1#7(A����sf|J7����YI���ϵ��~on�>��P9��$-1^͜r=u�2�.a8ǌ�#�fC���0�o-�הXe�	�+3���'�@qP��'�9��,n���A�Vj"��ՕJ����"-yu<�ch|W�-��7�+�z�ڢ�����)�uC\��1��9̂�1W�?`��Q�lNS*�lA�>"�p~���'	���7�z�������~zL-b?���J�2z�b�"̸O񒘩|����Aw	���[7,�B�r7�>�Vb��3?�������S��� &��GT�F��deÙ-�(i`���*-�0�%+�g�M��j1�Bs�W�d�K���C�Ey����M� Y"��B#iU�T�_m�� �Q�%P�5����V�Z/
�IkZ�>�}{6k�z2���c�5�^7�D�xQ$�
�Vd���m � ���Hx�M��D��]��{������}��%u�'��(��$Ж�	4A�m���vt U�Q� `>/��zC)l-�G���D�S�I�.-��J�-QXg
5N8׃<�Pf�P"Q@�.}����2����9e�x�z�����Cg�z�F[�f�J��/���Nq��-Z{\�����0�c�>���h�w?�$Vv��8;\m}�`  4[vVa����8F}:���tv={ �l��C%aN�nEt��L*7�=����ݦ�܊�%�)�eʣ��4�#�&O��DF()%^�q�_P�1�rŬR��)Tq ��;���ȟ���ӷ�����+�)�����?z��s�*	N��b6��q�߰��2 ��&6���W~s�ѫ��<�! &���SK���ڋ�R�� �+}��Uq��O��*��im�5Z]I>Я�ՔK���RtqnF���\��nÞ)\��#�AF�f�r�b?E|C�<,�4+�Q��C�����L4ղ���o�yz����M����$Z��Qc�\�u��N1���!K	�mY~x@b9��W�he)i��IYɛ.��bxI&LΩ�G8UA�b�	�6P�%����/���07K��U_�a��~�o���#̲W���3�z(0r����x���Oc<���dc�Ie��B��B�ҐT#{L�1��R��R�J��f(Sŷ苰ucM�N���V�r@J.
A�$�[�G\pʶ��B�Qf��o�|av�)��&�\iթ	NZ�`|�U`uSAղϯ���Xb���B��N(�!�x����_�𘿘

�=��[E����]�0�wܪ�wn�ﻥ(�u�LN�2zABBp�"��
�L,���Θ�BNV��7��4�/�|�_m.w�	@8����1�=��f�����j�ju��e����&#�Y�u�y̅�F�Y���c���"��.�m������A"��Ǣ��e��	>8�Em,�� ��
��J����h�jbo��zZ����H���L��+����K8������/k��)��IhE(�������Q\=H�
���;I\�-���Re�ʠ�����i�!6��.J��=f;�+bෝ�7,@Ș�oM��2��lA�6�tFp�hLj^p����m����mry�fj��e�N�,H<��S��yσ�_'�#��^�dZ�J�ֹ�^5�q݂C��f�*�;/Fv�5cPm�S��y}虸y���j��ì�Y�����L�>e}g>�S���tS
-�]�G}���/C�\�ܯ���X���-��0GCw��1�����]������bN��ŝ_6hC��&{ux|�3�is[y�7\�8[k�n��L'π-����/��lu{N���Ͷ|!I �OOW�-Sx���(N�I9cV�[���{�_fF���ƣ"�o���3���)N�k�u��8�`��O-����b�se�-,Ǳ�8���lF�=�X����ó���\Z��*ݣLŏ��E$d־�<�Vf?\/oM����j���(�`SK�����-A�!y-��.���4èiĳϔ�_�TtT`6�gD�W��QXL���(®U�	V�))� /WQ	�f�m����f��Zܪ��)�״
�<R�+\Z�w5�VI!Y�I$:���~X�qj�i ��+������qPɊ<�Y����+���� F�>�ŀ��P4�'p��!j��F̭C��<i����"%�1��z��'��<S�P�y`���8�����`B�߾
�d�H ��}�hK��}����*|"�f�[��0$��9_, �R�h�6��%akg�$�V��{�� �t��	@<�S�c�p��ܻ�2*���.`���h������=!���M�s��U�F|�|�5F͵o�%F���O%�$وM�Hγ�CN%�:�y���O2%t���lW��ik"v�'����e���K��kV#�=E�d��;\��ͽ�N'�s؋�^C`"l�;��C�z�j�k<ES�$�-~��:�&��H'�¹��$
9�"tx��I�`b���L��S���î��_���ͦ��D�K�����ȍ�+x���r�����;�3��js��4�o��_��v��X�{��k�����vE*���vQ� lV T\j�$*�ڠ�'�8yG�/{��Spe��a\+�<�a����	~�څ\s"��7ә�Ǯ/��]-#�jL�!�Kn�k�