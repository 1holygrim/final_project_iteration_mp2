XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����,��ҧ��E�8\��@�7b�P
���FOΕ��*��&��� ��6����}�$�ߦ��e!sK�(��q����g\n�_[L�?Z <s��ٞ^]��;�GY��']﯈�=P�\���ęEX���U��8�����V��+)I���X��T���k�h���`��j���8W�~f3���є�]y����B�T�~��	���  �<ۓS��ɗ�t���Kǚ���d�!,ُH3����!����~f��fj9��kW��}��\�#��nR�5��ʐ�!���.��c�
tV��~���� u�l�*�mYJ�w���{}Lk�S�z�>�<����vF�/�Ά�:���~�^�C�CD�WQj
�Ϡ��m��v'�Q���z�b�R�k�k�y�,�z�be�ՆT�>#?�u͉b$��C���.�!���cnҧ�{��R%�������Ϭ��+�Iq�cO�VE\�����jg�m��JZ���7�fˢ��+0o�)��O�8�~��"n7H�x�\	�U�.����NƢcY���DD�lT"�m}EC�A�G����qy��5mnM�v�V��������YQ )����6<e("��*���V2N"l�*�.�=cuJI��L!���$9�|����w�Y�7G9u��cˑz�?�,�Ya�6���;�� ���v�\�VÎ�g0L�)u'��yOL&��!��FX�51u"����d�y?Iz!��#�*	�JԱ��Դ�B�߶GXlxVHYEB    fa00    2a40�M ��fZ���y�&}.G�7���a�T����&4����-|�|W���㏕ {�����)�V�5�ݜT��t	(�!��
\l��(K�Xiw�I���ɡ��%�O`�$�wFf:Ic�� i+�K���w?�T>i�x��?�ovJyEK�Ltά�4Z��5��>C�ȳ��8�u5w��P�;��#�Iv��|��z2��Q�$�'���@�$���ĄTiu9ϷL�&v��2�C�Y�|V�\��uF�:�*)b�qZB��F��ҳ�[�����2o2C�b��;g!�٣^h��}�#�-�@��7�/c��J�2�X�K��&#���<�b=����A J�=I�]-M�;����m��V]�+٣����PL+:�Yj�j�ƅ����yLqEO?@��;��]�`��[�s(�; �8cNd��_Oe����$�'��4�<������U�X��2ͻ"s�YRU2�W��Y�&Tw�m�� ��������EB�O����T�? ��$�A'����5��8d:���R�8?�Pm����0y�b����+��mJق*���o� ?~xK �&%����1������I4w\��`���u�(X[|;1qݽ�N����a���p����wdlg��U��7Zb�q�Y�I��x?��T�<��V���iʇ=cu��8��p�
���P^����3V(�re^V����YλT� �{�dnٯ&���p����ÇejM�ۆ(w����!d*J��(��=�.��r)]q�_����Pl�	��p����g��ǯ�D����H���]��X3�y;�s�����D"�ex�3�ˉ
혤a�S�I��PC��=Vʐ�(&�\w�Ov�*�m��$��F̻��uL��Ȅ�e�	&6b9#���;�N{�e�}Br�cO/2���TWqƞ����\)!e?���J�U�/٘g��p}�[�(5h:�bk/�'r��Y25�S	��T��2l�C�c?��1�ӾxVs*�� u�R����KY0V�'�N�ý��el!�*=��u�S���e� ���XV�Ef�	�a��q���iٴ��T�:Mv^���I�~2ڎ-kh\٧��v3̖���V��q�a����ϴ$rb��P�>�����+̢�j�R1[&*�=*��[	(ǃy�N�P��͸���vIO�%,��8�^�xN0��8&0�OHj2����m������!��x�*Â>2����#p8���v�+Hc�}�"�QV��X/��S�Z��

(����\���Ƚ��Hp�ů�.U�%;|B��חT��ވ���T2Z���nH(}'���cp�/�{�!t�A`(�5R��D���r5k�|���yu�+X�`U���f4*U�8(�J䖒��6�r��_(�s�M7���	��G��]9)�q�T�qO�����5���)���h	��DѱH^V�\�0�]����SG
`�ݒ0��>V b��ܹ،|?�n԰wQ x�;�B��W �������o8��hon�����:ᕌM+��������,I������Z�;^���@DYm
6G��Hnʉ�B��#�A�bŢ���3��G"��S2_�������q!:Z���J�G܁�w] Y�$�iL��ޥ	vK8\� 7������g��j��5�����V�:(�a�I��'��)K�Č��F�;0�*3��g�:�G#��N�jP�ӻee� y,ej�m���[!�?A���:e��z�Q��0��v��3�L�|��7$C��n�7�y��;*h(.zk�߄a��=Mٟ��o�Xr�t|M�o8=�����ܐ/�0��8�3����ao'�V��TLmj�0�����>�B��$��W�Y	i��Km��ye�^���R8����m� v���@��,R�ř���mq��CEH��2/�K��	����m@&��#>�ȋ�A>�LOAE�^�wnO�g}]��p��}���k'm�ܝA��>]�i�x6��2�g`�8<�i�O�Z�[ ����w�����t��Ջ��o���Q��"VL2� _����:��j*Ƶ�̞I�M�D�n�(��]�B�1,�)C�����(��W�,����">@���l�V�Z�x':��}6+v%� D��s�8�f��HO����R>��'�)���[͸$��o^��v�hk�5�[Bw'2D�*	��&y�ɨ7d!,��)޲�k���>ʠ����+E�M��/�L2�ì\�������ӭ���p7�2&��=��>eډ����a�?���p�n���H�9�U�.tf��'�k ��{���!�⾧͖z̉�|���ejLB*�����S��xi�&`�Oz?��P�'µ	�%���1<���w��3X��f<�A�����
ŨJ��w�&����G���A]��s�����l�7d���)o71�]�P��L})D�S�P�gs���K�,��~���ɘFf�4���#�1����hu~�����n<�~�	�k����ʔֲ�\�D�
ԁ�+k�R3���zI�lhҨ��� y�:
o� 0�y��PEi��
�~��K�/P+��ʍm��,
����12"K;L�񑚗�6j�	+e	�0<w#u�ӊl����p>���/D�h�JX��!_�c���
zj�[P�G�Y�H�p4Yãح�B|$�u�
��-u�b�cS8�����L�����[�JM6�HA����U�mc~r���s�j�Zc��~��NFP/�g��W�Q����Km\,�.��K��q���Z��3���������T��%�d%���5��n�:�<Z�W�f���z�/�B�rh�����SF[��a	���rm�iL��Fڬ����6��q�
�z��=�����p���,֞?E�"�����^��"���v&�
��_5F2&A�I�0��`�T�=�k��
e��.ǛW$l�E���C�Y������iwH&�� Vi]l���[Ƃ� މ,�� �$n��2�AহC���1AS��ɳ���迤��@"���6��*�ƺ�<9i�!���_D|7�8���e�졧����ğ��v����W��{v筠��?�%s,��y�!�O~���:�{�Nr�=Y�8�#.����dn����-bD�:ZBxKQ���ߜ��j�TH�#JA��\�=�~�+��7�(hF��t������êp1�K
#�Pq,�J=g�Im�A�0�h�\Xj��j�����Q�vh�	@��Mn1�
{-/��Sg�¤y�T)�2��Y���43߄�a}Y�\�@�&��}�*;M�����_*�	�Ł�d���PyY=��V3���ٍe��#�F9d+�G+���� 傤�i���k<?�n����A�+u�����f�W�yx���[b@���];.}�����hp�ǳC�&D�z��/q��P��.��E��Q.����g[x{��͢e1�;2��i�B��Jɸ���V��K�xl!5/��f��[%	m�u�t	�Ly޾3.x8MK� ��
�8�~�lVNʭ֋'�>�:PvȑG��BG�$ `��ߗg�M>��t|��h��VA`;.����2�a���b-w�H�lڥ�T���{�-��k��Ĭ?]NK|�]^\�jB�s�O��'��=X��~�lY��k�Idom�ʧuS�)����k[�`�2@�3����W�ۄBm�ԇ~�Q�E���)�fP�r��vJU��l|'����<$��{sF���w���ٱ�,���F<�#Ɯ"dF
�>�k�*��;d��
q�KWx�
f�ªh����hCX·�b����'��忡F�Q�CI���9G��M+'��ρ�����w%��d?(����:�,�\�� S`�z��b�c�B�z��u}30:ї4�&k��҄P��Tu��qrR���O^�4�Q^�f|qK�
�Q����"�J�2�#���Ae��v��{D�᳖Ԛ��}�aIG�G��������se_<G ǖ���\�5���>@t���h�[?�H�;ǖ)�>��^�&f������T��c��mu�69SA��H�lm[Sk��ja�5J �� �ի��mkۂ�����f�j���&��M�Q�=���	,kI��Ϣ��3ߡF�0dh�r�tKS��ς;/R	K�t���`T.]?��-��\��Y�'N�!���z���-����Ӏ���}�[F�z��8���������g�,��QK�<�=-��v�y��k��R�ZTX%/��O��Z?-�4�y�D��h����,5Jv8�v:O��1 1���[t�r���8d��e�����qַ�I-���c=,��ʏ!��cpD�a0]قʢ>N�z�l�H)����H����*�h��V�3x�q��ER�� ��J��ޖԗ�{TV�c텈�^�����0��	�X��*qus`���l")��'�0��"HJXC�<� ��g?�!��nK�x������k��^���L�N���S��f�zy]��8����ZJЂ�x�f!)?:��a�����y	1{��1B���<>쥟�,JY�y*���u��`sV�n7n._�m�Æ��|��y[�]+e��d���1����S_�G*��o�̑���9 y���D�jU�X�2<�`�/K2aFf�+˶�
#V��0S�C��c�� ��	�fҋH6�{[Z�B9r�n��Ä�--EtB&�+$��3�
փ���=�Dj'�х-�"c�k�xp'��[A�Ǹo���q���n������0��i����@���#�#ȷ!��(��`������X���-�u���
���c����Y��w���N��;����G/ֽ�f=����M����1^Y溦魥����%}�RN0q�J�A�o+fH�����v�@�����\�n�WQ�j�T�r0�+�3�Yj�.a�ߊ���l=�����Y+-X"��Ʉ��}r1C)�Z�����d���B�]��)Ӿ��Ҥ� ~�b$��`w���}2H�����06�bZ\��Q�(g�v��bXb�y��C�{ŲpL5�w�[���q®��N�׼W���̥f����wH~c$[ĊF��� c��}kOE~G'Є��$<p�3��4| �H�3Z��G�M�]X�B[��
"�o^�u��rc���5��,�6���bf
����7�$6���q]�������� 6	�5(�1Ǜ��7�ʟh�f�x�����XК�hwa��0x?���.���B%��6s�J��l�S.��W�C�7���PBM0��sX*�^�P���^Gr����g��s��;M�..�X�Kn�G�P��>�}��Z�>�γ�^4���T9��������Y����{�#�����bzmj4C�)ԭ眃���	�L;�ܠ�M��;މ����٧]L�f�1 }�Q`E\k°�K��v�N��o>		���!v%SSK�)�b9��3�WI���ޒϸ��>�≫�`��P���;c��^����̂��X�`��j�{�q�U��'���K0�`���8��Y�Z)�(����jRBM��ۼ�p;�꘭�����j]�/�.O:8�i��}���k;�����έ?��aw��� �H=�S\�@���`S�WULAQT��x�pZ�6��0�G�D��z�!	<�V�)R�=�;�@��"v����&�z��6�)S�"���^//�Y�YaW�W9���k:;����<Z5�ѾT?���t�ʒ
�B�����2#n�6A��O�CGW�?pʋR��e�_0?X1`��s9z��A�U�47_�׎��^d�}�6����v6�o����ӃK%�Ղ�qT$lӹw�.n�/c(8ğq��eb�H�(]����I�6I�OK�,a���_���㇯�����cP���V,�f^QKL��0�0&�U����&�f�-��Z}rrUl��o�(��-9�2��`���4���q��VϽ[���~	:���Z��=z���x�;Np�jg��LKu���/��T �E!�g�Q���Ef���G�C�'��l��"G&8A 6��C:Z$NA�zsx���Т1ޚ�1p����`���e)�Y�! t� ��ô[D���'|�ޯL�r^���oS���7lD����W�:J�4�vBbzȶ���MKLV�K���<&�2��k,V�E����S�ۃ8�pYC�d')/�MM+��o,�gwM�3���] �^��6��혛wUk�1���W�'V~��oi
m���4���@�O�ٹC\�T-�s��c���,�Dٷ�F������������Q"|������>V+�uv�6�A�)
(Փ9/�88E/3'1�6�u��BI������°�"@+~�٪T՟X��"�jf$�������,*�ka9����b���*��n#��>R���/�Tlߌ~uB�p��ZK�0'�S��k�S���!n>���sZ�U�K�ׅ��u��7��VQ��BE$�N�"��ĩ���3Dτ�ےj#�����l-�����ݵR	4�(`�RY��+��۳1�[7VbP'7H�6P��=��ի�9g�P]ٌP��;����}-;��#غ���򁍎�>}�ų���
K�ˆ�ゝ�����k��i��8M�W�S7��F;E�xr�̗�]i����$�n�"����m��QQTmr��2�Y��ǅ���2����&/�ݤ��=�*��v/Sp��^�u
���(�::�t^���O2��_�������C*)jk��~��	ZTp�I��Z�!r%��A:T��=/Ʋ�Pm (z�">%��hE|et�4O{�t%'֦�����Fάg|�q[χݏN�]xcd��]"6�M*fZ��>yK�c�4�nw
�I���^�����Y$�f��xZb���SP�}�َ{�ܙ3j~v\��{�!��;�C�(_w����L�چ81����[�:�[��YxY����~��nw	��`'��ֶ��~�V��gF(MX��Eow_j�2�:`-Ȧק��F��)��5B[��j4�Hυ�����a�+#��� &������g�y�tn��\)�������qQ�j�ά�0ʩ���z�;j�C�sP�ת�p�r]�����̎P��_�T�C�<�%�7���2n^���d�_��*��L�a����QY�ˋqJU>��I[k5�Dj�C�z�.[����lp�XY�x��.��
hL|]Ԯ"��2�SVIE�W�<Jr��@p��I �>����"+��(Ę�D!�ybs��~��f���BO���~=�Њ�z jZoif|�z�?���g�D����N�k�'����mjJ�Xb������!�l�P5u�T�5��S�$��acd�XAUr���� �Ӽ9�=��_!s�0
@���|C7�^]Z�{�1�xx�];��/N�	�2�rGha��|�R��Jb���<Z(�&��R�ES���z��.8�%o��؃�mDyI�@5B�ջ'�#n6?�Dl��T�H��Pl�*�x��]���e�.���ϳ�oRRwտ��>`���Aʏ�:�#b6�8RƑ�nǯ2Sg��`���x�c�g.��
���=�-	�R����w�V�����fF	g�����p��E�N�B��^c�-��C��\E�����t����BP�P����¦�h�V�.PS�4���Ѱ�$��c/�Kw���IǼ����';�����l�j�^Ǹ�3��O��S25?68���WU�T`�Φ��0^������M�M��<ŦZO�rE��m�iOS�����I�Uu��0��'�]�#'�0����G�(��Oa�Y�C�fd���T�EhQ�L������)���[�M���c}��l\T^�,Ű)2���9"�t{?��)F��\�\9-�g X�T0=z3܋��Hl�2j�1�v�S�4s��7�N�)���>#h�������}�r0�����|�P1mٲ�|�MEp[��D�r���$L�3�k���4x�ɸ��=�� ��O����n\��4m�!�&"�0�y
�rR��Y0u�#��k�zl�]&���!�o*k&VH�g�mO,<���6��� �>��~�g��O�'���ֳ��ӥt��!.غ�F�.�A�Tŷ�t�U�xL(�?nda���빤�������N���9&��͋�M����c�`��'���W��gН5�:�R&��6�WD�%���������K�G��W:�"�E6�K���V۸���8H��0��|CԛsEQ�L��ㄢǗ"�h��9��m(W;�8���}��*V�u��WH	w!���J*���ܕ�l�2f[-I/%���3�5]������k� 8�S^��M�I���]s�W���{�L�\���*����9_S6K���X:C����uzdpۨ^nZ;�O��6݂�� �%.^� �[ ��r�G���}�)f����Jd�����j�8��ƹ��_��7��z�*g(&v��Zv� ��eל����"��B@~���� 0W�k�|�en> ��瑑8՚}����Տ�{{�ht��q摘�0���-�~�\�z-$?
�ܻ�g����c�|�2��u���1��z[��";F����nc������Z&Jww�p��E{탁�dt0�WW��ȴ���w����m.H��q�E�$��J��f�o��Բ�S[�H)�VG|.���PQ�yi�K4�9|F�OZ���G�Vq���>�x��6h�b�Qn�[�M�v����O�⯲� �Y����^J=���;�{C�	�������p���?����E"G�1��l�ۭU���6���c�A	f�l��"کq4�
�9 .?�7�����F��9Ņ@�Y�1��+��unV|���}�?ZkRˌf����bH@�iD�]�fT6�(h_G�V�;��
}c}���4c��p���-��:��-+�)UE��;��	2wBM�WHk&�;�
�F��i���u�;[�a�j�Ow�"�_11��V~��0��O?��l�pU�^U����{z��ֈ�E�y<��9�ټN#��iy+��Ú��2Z�>R��@f�3Ѵ����P-���h��y��TݾlC� ���6P�~Jq�`:uoL5ܽ%EY�<�Ń��>°3��6%�'�Tf�mԎr%Wr��:ٮ["�v�G�����Tk��>��:������v�rp��55X�Fe�H���8��P�/#7�� ��'>���;�N� 1��������TQ����!M���[�,3y[���}��Y�ȟ%`u�BP������	��k�aL��M�v���3M��z������~�	&�
�q\��dQ�8%ɻ�5�te-dw��Ú�}����N�2rԕkƨ��� ��2���]5~�3۞�tj5���9��؀�"���y4e��)��QޢQ`�4L����JA¦)�\�Y������2M- �wft!c���Mj.�-I������3\u�_�-��|�y�V�.Oy�{�9J��6<��O��+N���g�@F�a1r!������,�����v���x(��#�8B<; ]���
��� $����,�h tY
D�$>���""g�%J�I�K�91G6i����A���qt+򅌆�11h���T%��	�p��!��Tn$�)z�[���N0�2ދ>�j�k%��Z�s�v �
�@
gm�5��ekKv���!���DB�����:B�IX�.�;^,"�����k��x����A�JsU3=�_M�U�8�*N���u����1��,�*3�%��	��T�)n
�DI�Q�w�,��_�6��;��ٿ<���p���r�
!P�vx�L�ŕ���{�e�{�kS���?'��9�{�4���i+���b�#G!���1s�lE��	��pTۖq�����K�Ϛ�I�u���X貃�$�W�L貟����m�$5���1�x0��b[������.t��u�Z]����o���T���ZF��rk�v BUI��|��7���q4��G�b*�5D%;�Avc"3��O��#<��f�T�����_��SʹQ����y������	��`��d�g���r��^���� ���KR����{#�F��Dq��w��D ����x�g�L��TeU�m��|�a�_>�@�2���S�'����?f#�q�ǀs.��%uV��˨��,l����r#�j��,9�p�fv�1W���I�S�ŝM�%:�ҹ�]�_c*���^@)�Om��L�*�����O�)$�x
 ��.vo�h�&w08Ӑ϶��e;��_��ײ�XQuuV��q�5��Y�_XB�p��Gm������h�������s�(.�n��k�G�;�=�l:�
l�<���j]��<vD�k�<��,'�!T�vٰcT��߬Z�(Uo����o^a��%�_v�޸��[a�>e"�~�d�_��"��=a&i��>�w�ޓ�.��k�~m��MYT�K���ZK�N�OF��Dd���	�Z�ٛ�AsN=��6҃���>B"�j���0�G#E���=����<Ն�s�*8g>ۜ�>�]�s

w`V'9���.R��C
�)�|��h9���y_���IA�s��mXlxVHYEB    fa00     8e0 �桙�Rn\���K?�e���9��?� nt�q���dHK� e�)�}�Q��"�k�B��dzٽ)��հ�և�����~a5�0)h�䱖t�¾�`A�T�������3��-NJ��k��a�� W�*�;o���䍸�e(�N�
m��`���/!��LP:e�q�Q��	-���Z>�������A�)�ae��~��`�2�b~��#��պ�ڳ�a�_�;a�&��0�,��ڌ)�b:;@É"~�՚����I�c�H/���O��b��O��qO���qg�����O\�)6��\O�n~z���|ET���g�3nw+4X�;X��h�=��^./;X��,���њ�.�ܝ>^8�����7G2
;^�emArŊCܘ���<8�qD#���}Q��I��*G�Ǣ���%���o�'\��^���1�!&�#�w8���ՏP8*�]�E&v���7�_<�f�A�%R'�mJv�`�P�G����2�D�Afu=�Y��`���J�����\�R	F|Fte��P;����R�[�8C�R�,0��V�b��S��ր�-kM�J����b� �W�ox0����	����?2������ot��k*wv�3$Bmz	Q�7�8[���J�"Ax�����:�m�q���]�#�_A)���g|�n��B]��'ʧmu��S��0��njZe�	���"����D���L.�����n�bu�-��P^�r> �Z��a1�KE��.�#J���S^����z�j7���ִ�7�2J
V�r1�Ց=}5:y~�v�rlc��j�R�S�N�ئ�����3��~J�4��ř��f{;��,���US��
�h�/LD<6w�艮Hf�#��X~oe���/��#��8;;�� �W+�k�IKN�@����d*=���
5�L��Ԏ��K�����,�r�[��w�'6�M!�>�%���H�eJ���BWPS��Req��k�f�����k�C��Ř�,��MW�m������Uɒl��Cn��6��F@�=�,PC7O\��)g���Yߜ@�I��P��,�|�^���.�hfe�Hd�Q(��?��49�i0]�}Ñ�P���	&�����U���X�5%vD٣Htʠ�\w�C&t	��n[N|�U�����P"cDϝ�;�����U��h�D�G��`̾��9u"�x�����l�_����x���Ɵ9�����-pEw��]u.�%��I��ʸ��M��T��M�<���6��x��s;���b��TDG��M�NXo��t���4����o�������H*߮V�V���v�C���^�44�?0R��@�>D���夽c�z,)�n�N2��
�æJ~��w�o% ):�??�����-Y� u����Ӎ�b��aF��l>3~�����73z���n��Wº����⿭��pY� Ǯ��_o6\�^��5q|���$'6�� ;D�	�����\j9x}^佟/\gj�J�n+2��}���坋?�vQT���q�րpla�rv^Go�ɜ\u�F��Ɇ�Β����I���	鹲 ���� �q
��ӹ�Sݬ�*��c��s>Տ:�ӻ���䦹�6����������p�w��~�&Z�F�v�	�Tus����NQ�-U;w���uz)
�l�l�@e�wP�L´ u�)�Y��*e��'~{�Xu۩;E\k�Y+�{�A��g͢yﻛ$�����af^�D2�})A�"j����a����"L�v��
S>�|���צǂo�v5L�1���7L�)���qC0�d���Fw�Eg�'�Pڷh�L��"G�0�+P�d��l�W�ی0l�%��������N���c7�&���-M����+��H����R���cv+���~c��O+M���G���R;Q�.@.�_<Z��8[�K����)f�,��w�1f���L������2��ًR��q7� ��S�%�H&?+l�~�%yS"Ir_#�k��L^�������v	�Z��G�UkM�������ॺ�|,���8���I~d&�Q�Q���B<��<E�+qr^��H?)4��҈W�J��;�ػ���ָ�����w�5���H�Aӊ�+x�����|v�X����Fm��[I魲��DBVT���q)���}44�5�{'�L�կŃ}�L�b���6�0�� /m�"R&��^u��;�6����HLpXlxVHYEB    fa00    1110dX�{p&;���-f��rh�!�t�#N����t�2��*��f��ܝ���^���R�v٠j�˖5���Q������y� ms��D�ȉ^��Z�	1��؃"��?FF���������k���A̋���fR����p�ղv�	���Ae�o�@�li�~־�[h�5mp
��C��|W�Le��;S��`��5��o��x(#�F�b%
�ZLW�(B������XL+%�wx���	yJ�O
�U�h	-�n���J�'t5	�����chJq!5H�v��<R �f�5 ������Y� Xk � o�ӵ'� ����z}�F�����z��^*M���V���h���C����W��+E�"����E�3��2�=�_p�Z�3���#�w�A�ʿ��Is�*����v����2� <�����V�6s���	w�Q)-��a�%���_���q�Q@t�L����X�H��S�tEvo1�Yu���,��ƺ��4�PJ�D�f��$�xI{��F�lI�P��N�������u$%&툊�)�gp�2���d����#T�5�b���{hB��z�y�ث7U���z��\�OEjH��;?��ͦ�0���H@hD��H�W�fT���%(�b��FF�{[ĩt�����|�b�q'/�Km�x��T��"���)x��*���<����6vy��-:�1��s����ʧ�-A�'��G�1K����+�o5\��y�(�J�c���-�������b��>Ia]�f��8�����X㚿�pTRŅ|A[%T�*��iB�T�_�M��`����H4\����~�')x��u���L��n.t�	���XE0��@��U�~�urp��Mg�9ד��Zx��?��������Moy��ET����2F	&E�p����D ��;�Ϟp�a���UC�`��㹸4�yT��(xN��Mz-��L��ۢ?�']��a0��7�����Ο2Z�2�T��^1Kv������k�����1�=�Y��QUs�ͻA�Y�v
���s�F���z/�x�+VZ�+�z��@`���-�]S��gd��y� '�c���w�`I8?qT����R=��������b��L��{qXfg����E��޷�$C9�W8]��'A$f�g���g$���2��u^�vW&��Q!A;�5;���AlV夾��{�ȗy8��kzv�>so���|Cu��4�Q��(�<��e��9 *0�|͒NXe�@|�!�a�7�kEg�{v ���j��,/Q���r��+�-�������&4J���,�]^�N���7�j���:v1 ��A��,!*^Z�?����Eu�
�������'�l�����g��~�N�i�ޫ��a�_��7������%Z���
��Υ���An�"	I�ZG�7d^�'}���B����t�n<�;~${�����<��r&�����g�6Xe��GE_n{�E��V:#|�I%)��1'Jk����:�F���f qD�d7�oMT]¾dK��S� ����ո��^��w������!_Ne ����R�L&�3C��긊$�PWG����/���9�M��Y��帪#�[/��1׏xa��V5�����0Ui �fg�O�4�/�rX<2�z�5�i���"�ZTB<vP��_q�'����T9�}������O��K��o<�}L�0�c��W-��7Ai�]�����g��K�(�6���v�U|�(:�Ò��N&�8_3�)!��a$�ͼ�O�v�;cXR`l[V,�"�N,`��)��ꚑ���_�/�����$���؈h��>�~�$bgI��
x����V�c�2����Yo�v��^Z��g5؎X�*s�#-�Ik��)G�qS�n�fDw}��޽�>!�&�{g�IJY��}'�Ԛ-��O��KQ���XlF
X�Do���z�3�u��,�~����UG$Sn�ͻ�򭴎AI7^(	Q)c�8�S���;,���7>ۡ�Xc�C���R��c�%�s���ӏ�)��]�P\�릀���r_
��=�ZǢb`��Nߟ䵒o�3<���?dF�}	��oRt���l�m��6׼~^���4Z��J��<�~�/TNU����"c�Z}U�;��~bK��x,�|�O��E]"�|#c�-��)?� �����/ŹGD#m�<��{IY����Tb�ðx*�@Ld������دszu���o*	:��9Eu+���=^o8r�Ԕ�l�f��â+W�����4BC9�0�~�6��4��O��'�d���`�m���H-V�m��X��{��8y��r靍߰{J̢�M���e���i���qr��Z)�;��1d���)m����'b� bf�ٰ�^C�Ku�O�¼�,5�G������6>mP�V���DuY�T��n�SBC��҆E˓,��P����T��R�!�����<}��r �ط�\���h�Vn��Zi}ӈ�1���p!^ �O�������4�K]�-�sӟd�ku�:A��^�?�����lQy s�!�vD|j��l�5[^�|��Q"�E�k�
�u���߳�����o��=^\T<f�4�$hC���9V��B��_ L�G0h�.V�!+�*L{�ڎZ�VS+g�I��V�+~�\��R�x}چ��zKΤn�����!�\�^{^?���a��ن���2>؎dV��3C˞�0��#\�* �G��Y�6���8w9F"�sG8�y�wx/�s����P��IH���|��G�{���r�P��{F��o���B�Ve,��׶5Ύ.�[�]�jH�O�ّ3j.�@,�`0�Lލ��WΈ�[_�6�֦F�ǝ�L�]�dUv4("�Bϲk�C��K��
�]�����f�ʮ���Lۃ�w>�۰�,� c�zKdg��7PQ�*��7�v�۲&1��j��D�ɥ�dW�Y~NIZ�^&q9޳}��\M>�o9���AOrTn��ŗ�E�����&v>��	��B�\�D8��EYJ�o�q�^P�Ѣ&#L�ds��Q��.��2l�Vj߫z��p��AG��]�J5���k+}��.~:��@�1��LfVQz{�+�z���5��ƅv�	��K3I[�
�LE)�\(����w4�>�OΈX��UB��r�ذ���p�^-��q�jp�.�-�.hMm˖(¶��R���b���3D�L�)_98g�b*I��F��ݠ�I�6���BW0�\]w��Ͻ��raU$��dAZ!,*�}[b��8��n?�-�dO*6����ܴ`v�#ӱp�D���,�������?i�i��	m�Nl�FSϗ���+��#W�b�4ܾ��V�胰��g��V�W�jz�48b��)��0�����xP���+�R���f/�K���wj�j��>��d��;�i�[�#1��#@pP��9ݟ�����v4_E^M0ʨb��2��I;'���@!
��u�d�!��
D�Pg�$�Ԑ�aCez8&�
-�͙ţs�{�����R�$6�7u9�>��hK,��4y������ى��+/�Y,��Ꚉ��9�r(D��y��hM_C������`2�|r�^G9HK�y��`khlM���C��${q}ل!�dSb���N
�lI�6'v�;N�;�5����cνY�f�Cr���.�ihðSk�G��'���ڮӾ*&2��7X�a���ѿ�(��nI%�!��it���:||� Zs��
�+�}����m:�k]M�1Mω9�=$���4ɘ<�V�p<��f�rw�C5Kkr/���7�q�Q���"��59ʴn5����f_U���(��3�2��!��C�Kb���q~��[ZT�y��T3�1v�n1.5�/�HIuθ**q������ O7!F��0ħ��jV���J�(���%2Q�6���h�X�%�p�������X�rD�1��%��]���y8_ I�N�Q�?wڐ���O2E�c��)o2�l]"`�ȓ�|��>s���I��>B�8�^�8r�41kC�Hh�N�42�����l"c}�2%���VB7���V���3v�-1���5�`"��
į�0^p�]Ja��>27r�6�Z�?uxM�G�N���q�R�?D�we��%�2fu�W�`EV�U,{H10$�p�?M�H�"�ڄ=n�I�cNj�.Np[����k�C�E,VU<��X�p��{gl���<Ұ4�
�yi����o�M����%��,�o�������}���q�}p?TZx'�%$�'XlxVHYEB    fa00     ca0��3��,2K�����	�w
�<T�x��l8��\UH&���k�R �=v�9��fɱ!��u�r��IW�H�<]8�s��5�\� M��Xl<Nn� =��t�nM-�V����l��ۢ<bCɖ�n�d]΂��A	*�:|ek��I��H �2�Z��K�!�
X�Feۙ�j%Z������K�9_�������󓢠���r1�k����L�6TG���<Zl!J�}i�d���/�h���%')p�,s�Y;��C��Ph�=s�7�k .h�[��+W�_���E5C��%G��₺�1�������긠<�a�1�����T�����#�u��cL�����EHX^��wY�=u~,��QT��]~�B\��'��eّ��\�S����&�;����B*{#��������fx���]���2��z�T�01�H�n_`J��p��3�::�)�Npa����ԩe��y%��4X�>�a�4�گO�ߪ������Oȡ?8�E.�a�;,����t��n�����ɋ���"h�l���	ܒ�\�	��UJ
�J�Yau����wbw��\��%�Saf�SȮ2-rFo
x��Y6���y�\TV�~)^&>�`	�|�q�%f&}�@�57�(��Qq�93Y�?���V�flGV/5hv��7
����[�"GL���z�0w~Y��c�7�z��Fe��u ��$�*�q^���;6|J��I�%h�.I�
�O�la;�@�"�}Z�I�	��u(:�# �q��1㼚ȹE�NW��`KncLt��9�?eE���(�>"�#�rNӮ�沩=-1V�C��t�<#�����x�d44�&	?z�8�4p��WNûi�������"�������1�
ղ�Z<���:�/�ڔAP�+��Z�1���L.
�ը]C���ej��
n[�EJj��S�=�B➸���JWZ��	21�M���
Pn
A3m��*�8.�뙊��N�V� ���0���X�&�sj�.�l� w�"���К\���Ϫ��<H1J�M崇�tu�x�6ؘ���c4��
�`��U���G��D��$����@����(cp��C�m�;�u�$I�sUwp����INCPj�񇶘Y8�K$c�ḧMRRp���>���Ef�ޯm�����4m���J
p��Ql��Jm"�$����h��~�D���K�((#���]�Ky+E`�v֗��u*�r_=�:� ���h�'�&����ق�E��0��v�#�e�3�I�<I�Y��ƹ؞�*�/kx�7�Pz#	���RG��2p?�o���^Ø$K�Is�����m�70݌����dp���.��C���zT�2\�u��]�o�*������z�kk�Ɛ�*�: 3�95�<��E\�.r�y���Ý���c��&�<�۪������.:ԧ���j6L�M���`��|Cm��Z+
���Ł+�<f�ab����o����=��_(��]���rǖ/X?n6�E�&Љ���_7Ef���r4ϔE��1&9��?�����]ut��#����=�ͪ��$�^5)�eD�O?L$�`��v�j�XC&��v�9I���z�"�����(($�b���*����Qj#�
Ҳ鶐驘Á��ݥ ��-Ѝ_��I��(�o �g���,�y\>s[��@Z㎸1+O$Q�F�RVg!�*>�3�̔
�,�
.R���;��h=p���.9�^G�ۼ�'�/7B����ڇ�m6�SB\�;��c��P�'�k<N��m���w6U��[��Tn��6˲2��ݩ����U�Kf�'������E��Έm���dZ~���p��ͥ��*S�C OE�����c�� ��0�YLn��^G����� $�t�Ɩ#��KVan��¨8�53�7e�b�F}d��;�7�*��R\���a
����~ry�Mbt�R/��!F,�c��R���ݡ<2"�s�K�9
�%��C�;�* *q�����1��2�'��{���k���j5k����rKc�e��� �3"�*��:Xr�����E�����q�/>�D�+��"�Z3�ѝ���0jZΙ�+@b�kV�������o���	��r.y�S� ��b�TA^�g�`��O�g�j.|�������[����,���D�  (k��3%�o�t��a�\N��6g���Ip:�V�8�9��������~(��)r*$t���[](�u���9(ĔYJ�t�B(97xN��	[#Sn��ﾆ�2�'^=���-�ZQ~�Y~E�aߌ�-`��FA���ydE�����N��$O������l��6]�TfU!�!�SS�>#~�+N��՗���|����>3�M���Jn�96-eM�xh����k���JEBuw�i�!+J���.`=��p��
�S���9���M_o)��Q�Y3z<����s������h����OD����u�5�H�w.a�>��qN�,������� �9b��u��(��V$�KKt������\з�K�񝱵�(�"�P�#�P��F�m��e��	4�/�Y�ڴ�;��&d�M�1dr����S=o�8���)���B��F���w?4Ӽ�H��8��TG��-�gm>v+�#${�z�@D<�����ܲ&rC�:,���c�Y��Ճ�z������/\D�t��}$��	���KCK�L$�l�*��}o�`m�˯: ��2�K�\�"tNs$�TTv���n�$_�3Ra����Q�R��[�T�������\���v��hS�����R�"��@���p���#�ʢ��͖�);�S 1�`xMx꜈0E�?�т^ƿ|0P'U��-5�|�::0�:�mBg�f����.�z�p�{��
��5N��3)!0�X�*���,�Q�G�ye2�!GX�u�>o
?-�V0�{3?]'�ikPwZL.�ΐ�>�0����ǁ�}!Ϛv���4d��_����G��	�F(��8���b�u.��4p���l��W;s������s���G�(Ym.v����+��I��63�2~���q�MOn�7���3Cg[�:��30ͦ;t�^eoG0���[���9/��tzQ`h��!lj;��$�'��.��~����^F��GG���b��a���^#K�XlxVHYEB    fa00     3f0��y������hT��5��5^��{�^OҠ��<s7��&W���y��T����pO���X{jRT4/�fTMc؁�pYt�Fcz��: �����ZX��_������O��A��uuV੍+�R��1�'���}
N��nB9B�
��?���j�o��$'f�DCORl�K"����׍�(UA��3�*+���Z�@u��z��X��+�7��*��k%R�FN'/>��$��C+�����.�p0N��=Bm��o��c;��3Y�t[� 0t���`m���u�b��Yx�V�|��J5cw���Ź���!�������]1ώV0�i�7#O�\A���uUz��I�S�+I+�w�sp.a�I{�����f)t��Ɓ�#�b��C5��hH Z\�f�����W��C����{y�9ۧ�Z��|��cȇ&�S���e��2N(��M����,ۥ����f�
n������z�hP��}�+as��-���𙿚<@n��}KD ��^��b��xvv�����O���оU�uE.1�n�s�- ��+�h���rѡZ�}9~z:Bl:Ʒ�����*z��j�䗘���PS��⺰���T!�ǫ�ո�s���bǧP�<�@6�\���<�*� <���]}��e1�H�찣O�#Оd��P�r���V�՜?�>�CsUj"�6k�7���Ћ�{rg�I$ĵ��LӺ �����3�K���-B�� ɸ~����r��. �Ȃ#���-<JWWnں�ot����YK��'`�j��W�u(�)L8���η���}3{�C�h�����
����W=��Za\F�:1H?�O�NêS?�P�3�㼁����]�f9	����L�� ��>�:yQG�V.�� A����F5����6�w�5&A*���,����ڤj5�A�:��gN�+���J�o�>�����⾩w	��xO�d�N����Z�HU�8ҫ�+iE9��E�E(EUǜXlxVHYEB    8096     b20��[���=�)�	���������LjPC@8@�%�][������r��B����2��T�- �|���>��!�Z��c4�TۻM,¡F�F�+�_N(Rm�N������̴aC�=��a`�%O���O����#)���\J��~Eï�P����K�E��߅�)9W�S{u�jVhc�Kj�[�ǉ3�.rS��3�������d�-���g=�:ne(��d��oBp�@J�|���o6�9)���>�c`��/���y�"�u��i��P+!�0����9�B�Ƽ�dOp�z"�u~�Y?/?�h#řuX�s7�[����ȔD6�ueѦe7t�cS6�#�
������/���|l�[�^v�,�x	��N�ۆ���B��nj
+{�tv7ɤ�R<N=i�/��o�á��I|���/]o�A��N��w�P�%�$��k�S)˝PD*�Ǹ.��CD:Q���չP�gc*��vB�%hj�݋�3s3��W�J<������e�4�Շ�߹ ��X��=}+Y�/s��k��ReO�����c�;�B;h�:Fa������;�S-᳘6Ju/~w�ب�%�cJ�[e�;t� �Y	���[lR���ԊO#�����g���g�O�����_�>A��T	2��)�C��\���pY�6�IS���7a������2>�w���H���p�M�����������}b�{���P���S�)�Oy4S�)�@�ڤp�!�oފi����۾QfS��}���i��}����S(�*�Ĳ	{�����+�����jQ��<��up�m`z���r���I��7��.�-�$:Y�v(�����♏fǺ��6��`;���bg�;��2L��2/�U)ʭ�7��F��=L��$c�:�7G!Q��w����8�r�I�VK%�����n����Ƈ��4�NO&��;�nQQ�>zVT��7�X�M:L�� "���&�w=��ZO�ʠX�Z8�q$���Ș}'�Q�g�ǈ��:�M��㦴<FYa�a�:�ӂ΍�=�Jֻ�;])�)�s�y���$5����P#�}��r��V+t�L	g;�r�V�W�������h>�a�<	��b��,p͡G���H-�໬�,��+�g���(	F�S��X�@��Sj�ו�.�SUn"2?�� �N�(�`DZ]q��o0,�ie=k�e�~fx��=�毦
��8}F�V�{��"�l❼bB3e�`���W�(�_�����^�_t?�k`~�y׾	�c����븪��*��ȹm�E�9G���6�A�4���Bu5���p!��)ك����-k�� 9�u�$$B�u��^S�>�@�Nh�,�O�;�Q����~Z�߾T��Mi��!o�rf��w��Rγ{PBi�1�N���/_wR�]��T;��j*2_}��+HдT8d���[����¶�1i9��BJ��������"x���|�o�T�|Θ[�q���mH0ځÕZ�Di��qz�T-Z����$�	��ņ�"�
�fh��m�����n(�yƲ�D���Y;�ctѹ�T���Ӯ�t�Tmm_@��B�υ ����?���`��c�n4o�j��ѦL}!˛��/3�U>��>=sm�0�[������7��e���AS9j�!*�l�
�|λ<�epA��G/���]�;$�hx,BsAۣnS(g��R�)�
��$}G֐��`��4G6:�d���=�6�x��k[�p�)"�p߾4"9�+���c#��]�'�QM���.����ӳ���� D�Ql'�7��o��z�E�.J���}�@A:>_���4�Wy�0�/C/7Z��*�\xTWË�V�(gͤOZ+��ę�0�p�����Tվo��TLc!7� ��&7�ղ&���KK�.������oˉ��ovT�=��E��1r���>�
I^.K��Z�9�'M�x�h`���_U�L��H4<�.g��B ��+(�|�2��x�]���!ٿXf�$���X:N�Ph�L1��ƥ���zT�r+L��A�B١~��w��/�|�x���}�&iy�ދL�J�?TT�;�VT���/�Y`�k��=	V�@��=�/uVM�u>-^2���Y)��]��ϙ�v����8[rr�P�������E<#O2�Ǻ\c!Y�x���^���U �5�q�W��X]�7�95���n8������<��"aǖuYE��ӽ 0%��
ݑ���M�P�[�k.֜W���5E��7<a5����"�=(H������9hDuE&��7֕�������Щf��6��L����t���"Y��eb���Ozq��'zc5�$��&U�3�j0!9�*�L��:M*:��Q�d&
g�<������4���<�BZ��ۈ@�ڑW5|Vӿ���6℣2�0�lr�m9P�%�O�zxY�nN$SQ�`�Z<h�4VU��&�-�m� ̕�}[�n_o�Y��x
�L>S�B��g�Bd"��Q��R��O67�����w�ġ��;϶��l��9�J��6�e:3�Y�^�kO�2�:"ԝL��U�k4�n�m����i5�|.+��L�<W�˅�q�`/iTv"X8G*z5��B�S��ҞM?>Wq!�YY�+c-v(�6[�6vη82����6�b-�������$C��`���K�m@�^9�<)I��>��o�`vejQ�S=f�i��h�~B���~U+�s&���Ǯ����4,���f^�:Ȝ�y�$��LŰ�:�H��d��o���L�H9�&R�^�����hx\vR�cm+���vS�
��d6�A��